package Toplevel_Config is
	constant sysclk_frequency : integer := 80;
end package;
