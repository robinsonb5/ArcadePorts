
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity MiSTWrapper_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of MiSTWrapper_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"3b",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"29",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"38"),
    10 => (x"20",x"00",x"27",x"4f"),
    11 => (x"27",x"4e",x"00",x"00"),
    12 => (x"00",x"00",x"12",x"24"),
    13 => (x"87",x"fd",x"00",x"0f"),
    14 => (x"4f",x"87",x"fd",x"00"),
    15 => (x"c0",x"ff",x"1e",x"1e"),
    16 => (x"c4",x"48",x"69",x"49"),
    17 => (x"a6",x"c4",x"98",x"c0"),
    18 => (x"f4",x"02",x"6e",x"58"),
    19 => (x"79",x"66",x"c8",x"87"),
    20 => (x"87",x"c6",x"26",x"48"),
    21 => (x"4c",x"26",x"4d",x"26"),
    22 => (x"4f",x"26",x"4b",x"26"),
    23 => (x"5c",x"5b",x"5e",x"0e"),
    24 => (x"4c",x"66",x"cc",x"0e"),
    25 => (x"4a",x"14",x"4b",x"c0"),
    26 => (x"72",x"9a",x"ff",x"c3"),
    27 => (x"87",x"d5",x"02",x"9a"),
    28 => (x"1e",x"71",x"49",x"72"),
    29 => (x"c4",x"87",x"c5",x"ff"),
    30 => (x"14",x"83",x"c1",x"86"),
    31 => (x"9a",x"ff",x"c3",x"4a"),
    32 => (x"eb",x"05",x"9a",x"72"),
    33 => (x"ff",x"48",x"73",x"87"),
    34 => (x"5e",x"0e",x"87",x"cc"),
    35 => (x"0e",x"5d",x"5c",x"5b"),
    36 => (x"4b",x"c0",x"86",x"f0"),
    37 => (x"c0",x"48",x"a6",x"c4"),
    38 => (x"a6",x"e4",x"c0",x"78"),
    39 => (x"66",x"e0",x"c0",x"4c"),
    40 => (x"80",x"c1",x"48",x"49"),
    41 => (x"58",x"a6",x"e4",x"c0"),
    42 => (x"c0",x"fe",x"4a",x"11"),
    43 => (x"9a",x"72",x"ba",x"82"),
    44 => (x"87",x"d3",x"c4",x"02"),
    45 => (x"c3",x"02",x"66",x"c4"),
    46 => (x"a6",x"c4",x"87",x"e2"),
    47 => (x"72",x"78",x"c0",x"48"),
    48 => (x"aa",x"f0",x"c0",x"49"),
    49 => (x"87",x"f2",x"c2",x"02"),
    50 => (x"02",x"a9",x"e3",x"c1"),
    51 => (x"c1",x"87",x"f3",x"c2"),
    52 => (x"c0",x"02",x"a9",x"e4"),
    53 => (x"ec",x"c1",x"87",x"e1"),
    54 => (x"dd",x"c2",x"02",x"a9"),
    55 => (x"a9",x"f0",x"c1",x"87"),
    56 => (x"c1",x"87",x"d4",x"02"),
    57 => (x"c1",x"02",x"a9",x"f3"),
    58 => (x"f5",x"c1",x"87",x"fc"),
    59 => (x"87",x"c7",x"02",x"a9"),
    60 => (x"05",x"a9",x"f8",x"c1"),
    61 => (x"c4",x"87",x"dc",x"c2"),
    62 => (x"c4",x"49",x"74",x"84"),
    63 => (x"69",x"48",x"76",x"89"),
    64 => (x"c1",x"02",x"6e",x"78"),
    65 => (x"80",x"c8",x"87",x"d3"),
    66 => (x"a6",x"cc",x"78",x"c0"),
    67 => (x"6e",x"78",x"c0",x"48"),
    68 => (x"29",x"b7",x"dc",x"49"),
    69 => (x"9a",x"cf",x"4a",x"71"),
    70 => (x"30",x"c4",x"48",x"6e"),
    71 => (x"72",x"58",x"a6",x"c4"),
    72 => (x"87",x"c5",x"02",x"9a"),
    73 => (x"c1",x"48",x"a6",x"c8"),
    74 => (x"06",x"aa",x"c9",x"78"),
    75 => (x"f7",x"c0",x"87",x"c5"),
    76 => (x"c0",x"87",x"c3",x"82"),
    77 => (x"66",x"c8",x"82",x"f0"),
    78 => (x"72",x"87",x"c9",x"02"),
    79 => (x"87",x"fc",x"fb",x"1e"),
    80 => (x"83",x"c1",x"86",x"c4"),
    81 => (x"c1",x"48",x"66",x"cc"),
    82 => (x"58",x"a6",x"d0",x"80"),
    83 => (x"c8",x"48",x"66",x"cc"),
    84 => (x"fe",x"04",x"a8",x"b7"),
    85 => (x"d7",x"c1",x"87",x"f9"),
    86 => (x"1e",x"f0",x"c0",x"87"),
    87 => (x"c4",x"87",x"dd",x"fb"),
    88 => (x"c1",x"83",x"c1",x"86"),
    89 => (x"84",x"c4",x"87",x"ca"),
    90 => (x"89",x"c4",x"49",x"74"),
    91 => (x"eb",x"fb",x"1e",x"69"),
    92 => (x"70",x"86",x"c4",x"87"),
    93 => (x"c0",x"83",x"71",x"49"),
    94 => (x"a6",x"c4",x"87",x"f6"),
    95 => (x"c0",x"78",x"c1",x"48"),
    96 => (x"84",x"c4",x"87",x"ee"),
    97 => (x"89",x"c4",x"49",x"74"),
    98 => (x"ef",x"fa",x"1e",x"69"),
    99 => (x"c1",x"86",x"c4",x"87"),
   100 => (x"72",x"87",x"dd",x"83"),
   101 => (x"87",x"e4",x"fa",x"1e"),
   102 => (x"87",x"d4",x"86",x"c4"),
   103 => (x"05",x"aa",x"e5",x"c0"),
   104 => (x"a6",x"c4",x"87",x"c7"),
   105 => (x"c7",x"78",x"c1",x"48"),
   106 => (x"fa",x"1e",x"72",x"87"),
   107 => (x"86",x"c4",x"87",x"ce"),
   108 => (x"49",x"66",x"e0",x"c0"),
   109 => (x"c0",x"80",x"c1",x"48"),
   110 => (x"11",x"58",x"a6",x"e4"),
   111 => (x"82",x"c0",x"fe",x"4a"),
   112 => (x"05",x"9a",x"72",x"ba"),
   113 => (x"73",x"87",x"ed",x"fb"),
   114 => (x"26",x"8e",x"f0",x"48"),
   115 => (x"26",x"4c",x"26",x"4d"),
   116 => (x"0e",x"4f",x"26",x"4b"),
   117 => (x"86",x"e8",x"0e",x"5e"),
   118 => (x"c3",x"4a",x"d4",x"ff"),
   119 => (x"49",x"6a",x"7a",x"ff"),
   120 => (x"6a",x"7a",x"ff",x"c3"),
   121 => (x"c4",x"30",x"c8",x"48"),
   122 => (x"a6",x"c8",x"58",x"a6"),
   123 => (x"c3",x"b1",x"6e",x"59"),
   124 => (x"48",x"6a",x"7a",x"ff"),
   125 => (x"a6",x"cc",x"30",x"d0"),
   126 => (x"59",x"a6",x"d0",x"58"),
   127 => (x"c3",x"b1",x"66",x"c8"),
   128 => (x"48",x"6a",x"7a",x"ff"),
   129 => (x"a6",x"d4",x"30",x"d8"),
   130 => (x"59",x"a6",x"d8",x"58"),
   131 => (x"71",x"b1",x"66",x"d0"),
   132 => (x"c6",x"8e",x"e8",x"48"),
   133 => (x"26",x"4d",x"26",x"87"),
   134 => (x"26",x"4b",x"26",x"4c"),
   135 => (x"0e",x"5e",x"0e",x"4f"),
   136 => (x"d4",x"ff",x"86",x"f4"),
   137 => (x"7a",x"ff",x"c3",x"4a"),
   138 => (x"ff",x"c3",x"49",x"6a"),
   139 => (x"c8",x"48",x"71",x"7a"),
   140 => (x"58",x"a6",x"c4",x"30"),
   141 => (x"b1",x"6e",x"49",x"6a"),
   142 => (x"71",x"7a",x"ff",x"c3"),
   143 => (x"c8",x"30",x"c8",x"48"),
   144 => (x"49",x"6a",x"58",x"a6"),
   145 => (x"c3",x"b1",x"66",x"c4"),
   146 => (x"48",x"71",x"7a",x"ff"),
   147 => (x"a6",x"cc",x"30",x"c8"),
   148 => (x"c8",x"49",x"6a",x"58"),
   149 => (x"48",x"71",x"b1",x"66"),
   150 => (x"fe",x"fe",x"8e",x"f4"),
   151 => (x"5b",x"5e",x"0e",x"87"),
   152 => (x"d4",x"ff",x"0e",x"5c"),
   153 => (x"48",x"66",x"cc",x"4c"),
   154 => (x"70",x"98",x"ff",x"c3"),
   155 => (x"f4",x"cf",x"c1",x"7c"),
   156 => (x"87",x"c8",x"05",x"bf"),
   157 => (x"c9",x"48",x"66",x"d0"),
   158 => (x"58",x"a6",x"d4",x"30"),
   159 => (x"d8",x"49",x"66",x"d0"),
   160 => (x"c3",x"48",x"71",x"29"),
   161 => (x"7c",x"70",x"98",x"ff"),
   162 => (x"d0",x"49",x"66",x"d0"),
   163 => (x"c3",x"48",x"71",x"29"),
   164 => (x"7c",x"70",x"98",x"ff"),
   165 => (x"c8",x"49",x"66",x"d0"),
   166 => (x"c3",x"48",x"71",x"29"),
   167 => (x"7c",x"70",x"98",x"ff"),
   168 => (x"c3",x"48",x"66",x"d0"),
   169 => (x"7c",x"70",x"98",x"ff"),
   170 => (x"d0",x"49",x"66",x"cc"),
   171 => (x"c3",x"48",x"71",x"29"),
   172 => (x"7c",x"70",x"98",x"ff"),
   173 => (x"f0",x"c9",x"4a",x"6c"),
   174 => (x"ff",x"c3",x"4b",x"ff"),
   175 => (x"87",x"d2",x"05",x"aa"),
   176 => (x"6c",x"7c",x"ff",x"c3"),
   177 => (x"73",x"8b",x"c1",x"4a"),
   178 => (x"87",x"c6",x"02",x"9b"),
   179 => (x"02",x"aa",x"ff",x"c3"),
   180 => (x"48",x"72",x"87",x"ee"),
   181 => (x"1e",x"87",x"c0",x"fd"),
   182 => (x"d4",x"ff",x"49",x"c0"),
   183 => (x"78",x"ff",x"c3",x"48"),
   184 => (x"c8",x"c3",x"81",x"c1"),
   185 => (x"f1",x"04",x"a9",x"b7"),
   186 => (x"87",x"ef",x"fc",x"87"),
   187 => (x"0e",x"5b",x"5e",x"0e"),
   188 => (x"f8",x"c4",x"87",x"e5"),
   189 => (x"1e",x"c0",x"4b",x"df"),
   190 => (x"c1",x"f0",x"ff",x"c0"),
   191 => (x"dc",x"fd",x"1e",x"f7"),
   192 => (x"c1",x"86",x"c8",x"87"),
   193 => (x"ea",x"c0",x"05",x"a8"),
   194 => (x"48",x"d4",x"ff",x"87"),
   195 => (x"c1",x"78",x"ff",x"c3"),
   196 => (x"c0",x"c0",x"c0",x"c0"),
   197 => (x"e1",x"c0",x"1e",x"c0"),
   198 => (x"1e",x"e9",x"c1",x"f0"),
   199 => (x"c8",x"87",x"fe",x"fc"),
   200 => (x"05",x"98",x"70",x"86"),
   201 => (x"d4",x"ff",x"87",x"ca"),
   202 => (x"78",x"ff",x"c3",x"48"),
   203 => (x"87",x"cd",x"48",x"c1"),
   204 => (x"c1",x"87",x"e4",x"fe"),
   205 => (x"05",x"9b",x"73",x"8b"),
   206 => (x"c0",x"87",x"fb",x"fe"),
   207 => (x"87",x"d9",x"fb",x"48"),
   208 => (x"0e",x"5b",x"5e",x"0e"),
   209 => (x"c3",x"48",x"d4",x"ff"),
   210 => (x"e5",x"c0",x"78",x"ff"),
   211 => (x"cb",x"f4",x"1e",x"ce"),
   212 => (x"d3",x"86",x"c4",x"87"),
   213 => (x"c0",x"1e",x"c0",x"4b"),
   214 => (x"c1",x"c1",x"f0",x"ff"),
   215 => (x"87",x"fd",x"fb",x"1e"),
   216 => (x"98",x"70",x"86",x"c8"),
   217 => (x"ff",x"87",x"ca",x"05"),
   218 => (x"ff",x"c3",x"48",x"d4"),
   219 => (x"cd",x"48",x"c1",x"78"),
   220 => (x"87",x"e3",x"fd",x"87"),
   221 => (x"9b",x"73",x"8b",x"c1"),
   222 => (x"87",x"d9",x"ff",x"05"),
   223 => (x"d8",x"fa",x"48",x"c0"),
   224 => (x"5b",x"5e",x"0e",x"87"),
   225 => (x"ff",x"0e",x"5d",x"5c"),
   226 => (x"ca",x"fd",x"4d",x"d4"),
   227 => (x"1e",x"ea",x"c6",x"87"),
   228 => (x"c1",x"f0",x"e1",x"c0"),
   229 => (x"c4",x"fb",x"1e",x"c8"),
   230 => (x"70",x"86",x"c8",x"87"),
   231 => (x"d2",x"1e",x"73",x"4b"),
   232 => (x"e5",x"f3",x"1e",x"cc"),
   233 => (x"c1",x"86",x"c8",x"87"),
   234 => (x"87",x"c8",x"02",x"ab"),
   235 => (x"c0",x"87",x"d1",x"fe"),
   236 => (x"87",x"d3",x"c2",x"48"),
   237 => (x"70",x"87",x"e6",x"f9"),
   238 => (x"ff",x"ff",x"cf",x"49"),
   239 => (x"a9",x"ea",x"c6",x"99"),
   240 => (x"fd",x"87",x"c8",x"02"),
   241 => (x"48",x"c0",x"87",x"fa"),
   242 => (x"c3",x"87",x"fc",x"c1"),
   243 => (x"f1",x"c0",x"7d",x"ff"),
   244 => (x"87",x"d8",x"fc",x"4c"),
   245 => (x"c1",x"02",x"98",x"70"),
   246 => (x"1e",x"c0",x"87",x"d2"),
   247 => (x"c1",x"f0",x"ff",x"c0"),
   248 => (x"f8",x"f9",x"1e",x"fa"),
   249 => (x"70",x"86",x"c8",x"87"),
   250 => (x"05",x"9b",x"73",x"4b"),
   251 => (x"73",x"87",x"f3",x"c0"),
   252 => (x"1e",x"ca",x"d1",x"1e"),
   253 => (x"c8",x"87",x"d3",x"f2"),
   254 => (x"7d",x"ff",x"c3",x"86"),
   255 => (x"1e",x"73",x"4b",x"6d"),
   256 => (x"f2",x"1e",x"d6",x"d1"),
   257 => (x"86",x"c8",x"87",x"c4"),
   258 => (x"7d",x"7d",x"ff",x"c3"),
   259 => (x"49",x"73",x"7d",x"7d"),
   260 => (x"71",x"99",x"c0",x"c1"),
   261 => (x"87",x"c5",x"02",x"99"),
   262 => (x"ea",x"c0",x"48",x"c1"),
   263 => (x"c0",x"48",x"c0",x"87"),
   264 => (x"1e",x"73",x"87",x"e5"),
   265 => (x"f1",x"1e",x"e4",x"d1"),
   266 => (x"86",x"c8",x"87",x"e0"),
   267 => (x"cc",x"05",x"ac",x"c2"),
   268 => (x"1e",x"f0",x"d1",x"87"),
   269 => (x"c4",x"87",x"d3",x"f1"),
   270 => (x"ca",x"48",x"c0",x"86"),
   271 => (x"74",x"8c",x"c1",x"87"),
   272 => (x"cc",x"fe",x"05",x"9c"),
   273 => (x"f7",x"48",x"c0",x"87"),
   274 => (x"4d",x"43",x"87",x"cb"),
   275 => (x"20",x"38",x"35",x"44"),
   276 => (x"20",x"0a",x"64",x"25"),
   277 => (x"4d",x"43",x"00",x"20"),
   278 => (x"5f",x"38",x"35",x"44"),
   279 => (x"64",x"25",x"20",x"32"),
   280 => (x"00",x"20",x"20",x"0a"),
   281 => (x"35",x"44",x"4d",x"43"),
   282 => (x"64",x"25",x"20",x"38"),
   283 => (x"00",x"20",x"20",x"0a"),
   284 => (x"43",x"48",x"44",x"53"),
   285 => (x"69",x"6e",x"49",x"20"),
   286 => (x"6c",x"61",x"69",x"74"),
   287 => (x"74",x"61",x"7a",x"69"),
   288 => (x"20",x"6e",x"6f",x"69"),
   289 => (x"6f",x"72",x"72",x"65"),
   290 => (x"00",x"0a",x"21",x"72"),
   291 => (x"5f",x"64",x"6d",x"63"),
   292 => (x"38",x"44",x"4d",x"43"),
   293 => (x"73",x"65",x"72",x"20"),
   294 => (x"73",x"6e",x"6f",x"70"),
   295 => (x"25",x"20",x"3a",x"65"),
   296 => (x"0e",x"00",x"0a",x"64"),
   297 => (x"5d",x"5c",x"5b",x"5e"),
   298 => (x"d0",x"ff",x"1e",x"0e"),
   299 => (x"c0",x"c0",x"c8",x"4d"),
   300 => (x"f4",x"cf",x"c1",x"4b"),
   301 => (x"d6",x"78",x"c1",x"48"),
   302 => (x"df",x"ee",x"1e",x"c9"),
   303 => (x"c7",x"86",x"c4",x"87"),
   304 => (x"73",x"48",x"6d",x"4c"),
   305 => (x"58",x"a6",x"c4",x"98"),
   306 => (x"cc",x"c0",x"02",x"6e"),
   307 => (x"73",x"48",x"6d",x"87"),
   308 => (x"58",x"a6",x"c4",x"98"),
   309 => (x"f4",x"ff",x"05",x"6e"),
   310 => (x"f7",x"7d",x"c2",x"87"),
   311 => (x"48",x"6d",x"87",x"f9"),
   312 => (x"a6",x"c4",x"98",x"73"),
   313 => (x"c0",x"02",x"6e",x"58"),
   314 => (x"48",x"6d",x"87",x"cc"),
   315 => (x"a6",x"c4",x"98",x"73"),
   316 => (x"ff",x"05",x"6e",x"58"),
   317 => (x"7d",x"c3",x"87",x"f4"),
   318 => (x"e5",x"c0",x"1e",x"c0"),
   319 => (x"1e",x"c0",x"c1",x"d0"),
   320 => (x"c8",x"87",x"da",x"f5"),
   321 => (x"05",x"a8",x"c1",x"86"),
   322 => (x"c1",x"87",x"c2",x"c0"),
   323 => (x"05",x"ac",x"c2",x"4c"),
   324 => (x"d6",x"87",x"cd",x"c0"),
   325 => (x"c3",x"ed",x"1e",x"c4"),
   326 => (x"c0",x"86",x"c4",x"87"),
   327 => (x"87",x"e0",x"c1",x"48"),
   328 => (x"9c",x"74",x"8c",x"c1"),
   329 => (x"87",x"d9",x"fe",x"05"),
   330 => (x"c1",x"87",x"d6",x"f9"),
   331 => (x"c1",x"58",x"f8",x"cf"),
   332 => (x"05",x"bf",x"f4",x"cf"),
   333 => (x"c1",x"87",x"cd",x"c0"),
   334 => (x"f0",x"ff",x"c0",x"1e"),
   335 => (x"f4",x"1e",x"d0",x"c1"),
   336 => (x"86",x"c8",x"87",x"db"),
   337 => (x"c3",x"48",x"d4",x"ff"),
   338 => (x"c5",x"ca",x"78",x"ff"),
   339 => (x"fc",x"cf",x"c1",x"87"),
   340 => (x"f8",x"cf",x"c1",x"58"),
   341 => (x"cd",x"d6",x"1e",x"bf"),
   342 => (x"87",x"ee",x"ec",x"1e"),
   343 => (x"48",x"6d",x"86",x"c8"),
   344 => (x"a6",x"c4",x"98",x"73"),
   345 => (x"c0",x"02",x"6e",x"58"),
   346 => (x"48",x"6d",x"87",x"cc"),
   347 => (x"a6",x"c4",x"98",x"73"),
   348 => (x"ff",x"05",x"6e",x"58"),
   349 => (x"7d",x"c2",x"87",x"f4"),
   350 => (x"c3",x"48",x"d4",x"ff"),
   351 => (x"48",x"c1",x"78",x"ff"),
   352 => (x"87",x"d1",x"f2",x"26"),
   353 => (x"52",x"52",x"45",x"49"),
   354 => (x"49",x"50",x"53",x"00"),
   355 => (x"20",x"44",x"53",x"00"),
   356 => (x"64",x"72",x"61",x"63"),
   357 => (x"7a",x"69",x"73",x"20"),
   358 => (x"73",x"69",x"20",x"65"),
   359 => (x"0a",x"64",x"25",x"20"),
   360 => (x"5b",x"5e",x"0e",x"00"),
   361 => (x"1e",x"0e",x"5d",x"5c"),
   362 => (x"ff",x"4c",x"ff",x"c3"),
   363 => (x"7b",x"74",x"4b",x"d4"),
   364 => (x"48",x"bf",x"d0",x"ff"),
   365 => (x"98",x"c0",x"c0",x"c8"),
   366 => (x"6e",x"58",x"a6",x"c4"),
   367 => (x"87",x"d0",x"c0",x"02"),
   368 => (x"48",x"bf",x"d0",x"ff"),
   369 => (x"98",x"c0",x"c0",x"c8"),
   370 => (x"6e",x"58",x"a6",x"c4"),
   371 => (x"87",x"f0",x"ff",x"05"),
   372 => (x"c4",x"48",x"d0",x"ff"),
   373 => (x"7b",x"74",x"78",x"c3"),
   374 => (x"c0",x"1e",x"66",x"d4"),
   375 => (x"d8",x"c1",x"f0",x"ff"),
   376 => (x"87",x"f9",x"f1",x"1e"),
   377 => (x"98",x"70",x"86",x"c8"),
   378 => (x"87",x"cd",x"c0",x"02"),
   379 => (x"e9",x"1e",x"c3",x"da"),
   380 => (x"86",x"c4",x"87",x"ea"),
   381 => (x"c6",x"c2",x"48",x"c1"),
   382 => (x"c3",x"7b",x"74",x"87"),
   383 => (x"4d",x"c0",x"7b",x"fe"),
   384 => (x"49",x"bf",x"66",x"d8"),
   385 => (x"b7",x"d8",x"4a",x"71"),
   386 => (x"74",x"48",x"72",x"2a"),
   387 => (x"71",x"7b",x"70",x"98"),
   388 => (x"2a",x"b7",x"d0",x"4a"),
   389 => (x"98",x"74",x"48",x"72"),
   390 => (x"4a",x"71",x"7b",x"70"),
   391 => (x"72",x"2a",x"b7",x"c8"),
   392 => (x"70",x"98",x"74",x"48"),
   393 => (x"74",x"48",x"71",x"7b"),
   394 => (x"d8",x"7b",x"70",x"98"),
   395 => (x"80",x"c4",x"48",x"66"),
   396 => (x"c1",x"58",x"a6",x"dc"),
   397 => (x"b7",x"c0",x"c2",x"85"),
   398 => (x"c3",x"ff",x"04",x"ad"),
   399 => (x"74",x"7b",x"74",x"87"),
   400 => (x"d8",x"7b",x"74",x"7b"),
   401 => (x"74",x"49",x"e0",x"da"),
   402 => (x"c0",x"05",x"6b",x"7b"),
   403 => (x"89",x"c1",x"87",x"c8"),
   404 => (x"ff",x"05",x"99",x"71"),
   405 => (x"7b",x"74",x"87",x"f1"),
   406 => (x"48",x"bf",x"d0",x"ff"),
   407 => (x"98",x"c0",x"c0",x"c8"),
   408 => (x"6e",x"58",x"a6",x"c4"),
   409 => (x"87",x"d0",x"c0",x"02"),
   410 => (x"48",x"bf",x"d0",x"ff"),
   411 => (x"98",x"c0",x"c0",x"c8"),
   412 => (x"6e",x"58",x"a6",x"c4"),
   413 => (x"87",x"f0",x"ff",x"05"),
   414 => (x"c2",x"48",x"d0",x"ff"),
   415 => (x"26",x"48",x"c0",x"78"),
   416 => (x"57",x"87",x"d2",x"ee"),
   417 => (x"65",x"74",x"69",x"72"),
   418 => (x"69",x"61",x"66",x"20"),
   419 => (x"0a",x"64",x"65",x"6c"),
   420 => (x"5b",x"5e",x"0e",x"00"),
   421 => (x"66",x"d0",x"0e",x"5c"),
   422 => (x"4b",x"66",x"cc",x"4c"),
   423 => (x"ee",x"c5",x"4a",x"c0"),
   424 => (x"ff",x"49",x"df",x"cd"),
   425 => (x"ff",x"c3",x"48",x"d4"),
   426 => (x"48",x"bf",x"70",x"78"),
   427 => (x"05",x"a8",x"fe",x"c3"),
   428 => (x"c1",x"87",x"d8",x"c1"),
   429 => (x"c0",x"48",x"f0",x"cf"),
   430 => (x"ac",x"b7",x"c4",x"78"),
   431 => (x"87",x"dc",x"c0",x"04"),
   432 => (x"70",x"87",x"d0",x"ec"),
   433 => (x"c4",x"7b",x"71",x"49"),
   434 => (x"f0",x"cf",x"c1",x"83"),
   435 => (x"80",x"71",x"48",x"bf"),
   436 => (x"58",x"f4",x"cf",x"c1"),
   437 => (x"ac",x"b7",x"8c",x"c4"),
   438 => (x"87",x"e4",x"ff",x"03"),
   439 => (x"06",x"ac",x"b7",x"c0"),
   440 => (x"ff",x"87",x"e5",x"c0"),
   441 => (x"ff",x"c3",x"48",x"d4"),
   442 => (x"49",x"bf",x"70",x"78"),
   443 => (x"c3",x"7b",x"97",x"71"),
   444 => (x"83",x"c1",x"98",x"ff"),
   445 => (x"bf",x"f0",x"cf",x"c1"),
   446 => (x"c1",x"80",x"71",x"48"),
   447 => (x"c1",x"58",x"f4",x"cf"),
   448 => (x"ac",x"b7",x"c0",x"8c"),
   449 => (x"87",x"db",x"ff",x"01"),
   450 => (x"c1",x"4a",x"49",x"c1"),
   451 => (x"05",x"99",x"71",x"89"),
   452 => (x"ff",x"87",x"d0",x"fe"),
   453 => (x"ff",x"c3",x"48",x"d4"),
   454 => (x"eb",x"48",x"72",x"78"),
   455 => (x"5e",x"0e",x"87",x"f9"),
   456 => (x"1e",x"0e",x"5c",x"5b"),
   457 => (x"4b",x"c0",x"c0",x"c8"),
   458 => (x"d4",x"ff",x"4c",x"c0"),
   459 => (x"78",x"ff",x"c3",x"48"),
   460 => (x"48",x"bf",x"d0",x"ff"),
   461 => (x"a6",x"c4",x"98",x"73"),
   462 => (x"c0",x"02",x"6e",x"58"),
   463 => (x"d0",x"ff",x"87",x"ce"),
   464 => (x"98",x"73",x"48",x"bf"),
   465 => (x"6e",x"58",x"a6",x"c4"),
   466 => (x"87",x"f2",x"ff",x"05"),
   467 => (x"c4",x"48",x"d0",x"ff"),
   468 => (x"d4",x"ff",x"78",x"c3"),
   469 => (x"78",x"ff",x"c3",x"48"),
   470 => (x"c0",x"1e",x"66",x"d0"),
   471 => (x"d1",x"c1",x"f0",x"ff"),
   472 => (x"87",x"f9",x"eb",x"1e"),
   473 => (x"49",x"70",x"86",x"c8"),
   474 => (x"c0",x"02",x"99",x"71"),
   475 => (x"1e",x"71",x"87",x"d0"),
   476 => (x"de",x"1e",x"66",x"d4"),
   477 => (x"d1",x"e4",x"1e",x"f2"),
   478 => (x"c0",x"86",x"cc",x"87"),
   479 => (x"c0",x"c8",x"87",x"ee"),
   480 => (x"1e",x"66",x"d8",x"1e"),
   481 => (x"c8",x"87",x"ca",x"fc"),
   482 => (x"ff",x"4c",x"70",x"86"),
   483 => (x"73",x"48",x"bf",x"d0"),
   484 => (x"58",x"a6",x"c4",x"98"),
   485 => (x"ce",x"c0",x"02",x"6e"),
   486 => (x"bf",x"d0",x"ff",x"87"),
   487 => (x"c4",x"98",x"73",x"48"),
   488 => (x"05",x"6e",x"58",x"a6"),
   489 => (x"ff",x"87",x"f2",x"ff"),
   490 => (x"78",x"c2",x"48",x"d0"),
   491 => (x"e9",x"26",x"48",x"74"),
   492 => (x"65",x"52",x"87",x"e5"),
   493 => (x"63",x"20",x"64",x"61"),
   494 => (x"61",x"6d",x"6d",x"6f"),
   495 => (x"66",x"20",x"64",x"6e"),
   496 => (x"65",x"6c",x"69",x"61"),
   497 => (x"74",x"61",x"20",x"64"),
   498 => (x"20",x"64",x"25",x"20"),
   499 => (x"29",x"64",x"25",x"28"),
   500 => (x"5e",x"0e",x"00",x"0a"),
   501 => (x"0e",x"5d",x"5c",x"5b"),
   502 => (x"c0",x"1e",x"c0",x"1e"),
   503 => (x"c9",x"c1",x"f0",x"ff"),
   504 => (x"87",x"f9",x"e9",x"1e"),
   505 => (x"1e",x"d2",x"86",x"c8"),
   506 => (x"1e",x"c2",x"d0",x"c1"),
   507 => (x"c8",x"87",x"e2",x"fa"),
   508 => (x"c1",x"4d",x"c0",x"86"),
   509 => (x"ad",x"b7",x"d2",x"85"),
   510 => (x"87",x"f7",x"ff",x"04"),
   511 => (x"97",x"c2",x"d0",x"c1"),
   512 => (x"c0",x"c3",x"49",x"bf"),
   513 => (x"a9",x"c0",x"c1",x"99"),
   514 => (x"87",x"e8",x"c0",x"05"),
   515 => (x"97",x"c9",x"d0",x"c1"),
   516 => (x"31",x"d0",x"49",x"bf"),
   517 => (x"97",x"ca",x"d0",x"c1"),
   518 => (x"32",x"c8",x"4a",x"bf"),
   519 => (x"d0",x"c1",x"b1",x"72"),
   520 => (x"4a",x"bf",x"97",x"cb"),
   521 => (x"ff",x"cf",x"b1",x"72"),
   522 => (x"71",x"99",x"ff",x"ff"),
   523 => (x"ca",x"85",x"c1",x"4d"),
   524 => (x"87",x"f0",x"c2",x"35"),
   525 => (x"97",x"cb",x"d0",x"c1"),
   526 => (x"33",x"c1",x"4b",x"bf"),
   527 => (x"d0",x"c1",x"9b",x"c6"),
   528 => (x"49",x"bf",x"97",x"cc"),
   529 => (x"71",x"29",x"b7",x"c7"),
   530 => (x"c7",x"d0",x"c1",x"b3"),
   531 => (x"71",x"49",x"bf",x"97"),
   532 => (x"c4",x"98",x"cf",x"48"),
   533 => (x"d0",x"c1",x"58",x"a6"),
   534 => (x"4c",x"bf",x"97",x"c8"),
   535 => (x"34",x"ca",x"9c",x"c3"),
   536 => (x"97",x"c9",x"d0",x"c1"),
   537 => (x"31",x"c2",x"49",x"bf"),
   538 => (x"d0",x"c1",x"b4",x"71"),
   539 => (x"49",x"bf",x"97",x"ca"),
   540 => (x"c6",x"99",x"c0",x"c3"),
   541 => (x"b4",x"71",x"29",x"b7"),
   542 => (x"66",x"c4",x"1e",x"74"),
   543 => (x"c0",x"1e",x"73",x"1e"),
   544 => (x"e0",x"1e",x"ea",x"e3"),
   545 => (x"86",x"d0",x"87",x"c4"),
   546 => (x"48",x"c1",x"83",x"c2"),
   547 => (x"4b",x"70",x"30",x"73"),
   548 => (x"e4",x"c0",x"1e",x"73"),
   549 => (x"df",x"ff",x"1e",x"d7"),
   550 => (x"86",x"c8",x"87",x"f0"),
   551 => (x"30",x"6e",x"48",x"c1"),
   552 => (x"74",x"58",x"a6",x"c4"),
   553 => (x"71",x"81",x"c1",x"49"),
   554 => (x"95",x"b7",x"73",x"4d"),
   555 => (x"1e",x"75",x"1e",x"6e"),
   556 => (x"1e",x"e0",x"e4",x"c0"),
   557 => (x"87",x"d2",x"df",x"ff"),
   558 => (x"48",x"6e",x"86",x"cc"),
   559 => (x"a8",x"b7",x"c0",x"c8"),
   560 => (x"87",x"d4",x"c0",x"06"),
   561 => (x"48",x"6e",x"35",x"c1"),
   562 => (x"c4",x"28",x"b7",x"c1"),
   563 => (x"48",x"6e",x"58",x"a6"),
   564 => (x"a8",x"b7",x"c0",x"c8"),
   565 => (x"87",x"ec",x"ff",x"01"),
   566 => (x"e4",x"c0",x"1e",x"75"),
   567 => (x"de",x"ff",x"1e",x"f6"),
   568 => (x"86",x"c8",x"87",x"e8"),
   569 => (x"e4",x"26",x"48",x"75"),
   570 => (x"5f",x"63",x"87",x"eb"),
   571 => (x"65",x"7a",x"69",x"73"),
   572 => (x"6c",x"75",x"6d",x"5f"),
   573 => (x"25",x"20",x"3a",x"74"),
   574 => (x"72",x"20",x"2c",x"64"),
   575 => (x"5f",x"64",x"61",x"65"),
   576 => (x"6c",x"5f",x"6c",x"62"),
   577 => (x"20",x"3a",x"6e",x"65"),
   578 => (x"20",x"2c",x"64",x"25"),
   579 => (x"7a",x"69",x"73",x"63"),
   580 => (x"25",x"20",x"3a",x"65"),
   581 => (x"4d",x"00",x"0a",x"64"),
   582 => (x"20",x"74",x"6c",x"75"),
   583 => (x"00",x"0a",x"64",x"25"),
   584 => (x"62",x"20",x"64",x"25"),
   585 => (x"6b",x"63",x"6f",x"6c"),
   586 => (x"66",x"6f",x"20",x"73"),
   587 => (x"7a",x"69",x"73",x"20"),
   588 => (x"64",x"25",x"20",x"65"),
   589 => (x"64",x"25",x"00",x"0a"),
   590 => (x"6f",x"6c",x"62",x"20"),
   591 => (x"20",x"73",x"6b",x"63"),
   592 => (x"35",x"20",x"66",x"6f"),
   593 => (x"62",x"20",x"32",x"31"),
   594 => (x"73",x"65",x"74",x"79"),
   595 => (x"4d",x"43",x"00",x"0a"),
   596 => (x"5e",x"0e",x"00",x"44"),
   597 => (x"4b",x"c0",x"0e",x"5b"),
   598 => (x"c0",x"48",x"66",x"d0"),
   599 => (x"c0",x"06",x"a8",x"b7"),
   600 => (x"66",x"c8",x"87",x"f6"),
   601 => (x"fe",x"4a",x"bf",x"97"),
   602 => (x"c8",x"ba",x"82",x"c0"),
   603 => (x"80",x"c1",x"48",x"66"),
   604 => (x"cc",x"58",x"a6",x"cc"),
   605 => (x"49",x"bf",x"97",x"66"),
   606 => (x"b9",x"81",x"c0",x"fe"),
   607 => (x"c1",x"48",x"66",x"cc"),
   608 => (x"58",x"a6",x"d0",x"80"),
   609 => (x"02",x"aa",x"b7",x"71"),
   610 => (x"48",x"c1",x"87",x"c4"),
   611 => (x"83",x"c1",x"87",x"cc"),
   612 => (x"ab",x"b7",x"66",x"d0"),
   613 => (x"87",x"ca",x"ff",x"04"),
   614 => (x"87",x"c4",x"48",x"c0"),
   615 => (x"4c",x"26",x"4d",x"26"),
   616 => (x"4f",x"26",x"4b",x"26"),
   617 => (x"5c",x"5b",x"5e",x"0e"),
   618 => (x"d8",x"c1",x"0e",x"5d"),
   619 => (x"78",x"c0",x"48",x"dc"),
   620 => (x"1e",x"fe",x"c0",x"c1"),
   621 => (x"87",x"e4",x"da",x"ff"),
   622 => (x"d0",x"c1",x"86",x"c4"),
   623 => (x"1e",x"c0",x"1e",x"d4"),
   624 => (x"c8",x"87",x"db",x"f5"),
   625 => (x"05",x"98",x"70",x"86"),
   626 => (x"fd",x"c0",x"87",x"cf"),
   627 => (x"da",x"ff",x"1e",x"ea"),
   628 => (x"86",x"c4",x"87",x"ca"),
   629 => (x"d6",x"cb",x"48",x"c0"),
   630 => (x"cb",x"c1",x"c1",x"87"),
   631 => (x"fb",x"d9",x"ff",x"1e"),
   632 => (x"c0",x"86",x"c4",x"87"),
   633 => (x"c8",x"d9",x"c1",x"4b"),
   634 => (x"c8",x"78",x"c1",x"48"),
   635 => (x"e2",x"c1",x"c1",x"1e"),
   636 => (x"ca",x"d1",x"c1",x"1e"),
   637 => (x"87",x"da",x"fd",x"1e"),
   638 => (x"98",x"70",x"86",x"cc"),
   639 => (x"c1",x"87",x"c6",x"05"),
   640 => (x"c0",x"48",x"c8",x"d9"),
   641 => (x"c1",x"1e",x"c8",x"78"),
   642 => (x"c1",x"1e",x"eb",x"c1"),
   643 => (x"fd",x"1e",x"e6",x"d1"),
   644 => (x"86",x"cc",x"87",x"c0"),
   645 => (x"c6",x"05",x"98",x"70"),
   646 => (x"c8",x"d9",x"c1",x"87"),
   647 => (x"c1",x"78",x"c0",x"48"),
   648 => (x"1e",x"bf",x"c8",x"d9"),
   649 => (x"1e",x"f4",x"c1",x"c1"),
   650 => (x"87",x"de",x"d9",x"ff"),
   651 => (x"d9",x"c1",x"86",x"c8"),
   652 => (x"c2",x"02",x"bf",x"c8"),
   653 => (x"d0",x"c1",x"87",x"d8"),
   654 => (x"d7",x"c1",x"4d",x"d4"),
   655 => (x"d8",x"c1",x"4c",x"d2"),
   656 => (x"49",x"bf",x"9f",x"d2"),
   657 => (x"d8",x"c1",x"1e",x"71"),
   658 => (x"d0",x"c1",x"49",x"d2"),
   659 => (x"1e",x"71",x"89",x"d4"),
   660 => (x"c0",x"c8",x"1e",x"d0"),
   661 => (x"dc",x"fe",x"c0",x"1e"),
   662 => (x"ed",x"d8",x"ff",x"1e"),
   663 => (x"74",x"86",x"d4",x"87"),
   664 => (x"69",x"81",x"c8",x"49"),
   665 => (x"d2",x"d8",x"c1",x"4b"),
   666 => (x"c5",x"49",x"bf",x"9f"),
   667 => (x"05",x"a9",x"ea",x"d6"),
   668 => (x"74",x"87",x"d0",x"c0"),
   669 => (x"69",x"81",x"c8",x"49"),
   670 => (x"87",x"d9",x"d9",x"1e"),
   671 => (x"4b",x"70",x"86",x"c4"),
   672 => (x"75",x"87",x"df",x"c0"),
   673 => (x"81",x"fe",x"c7",x"49"),
   674 => (x"ca",x"49",x"69",x"9f"),
   675 => (x"02",x"a9",x"d5",x"e9"),
   676 => (x"c0",x"87",x"cf",x"c0"),
   677 => (x"ff",x"1e",x"fe",x"fd"),
   678 => (x"c4",x"87",x"c1",x"d7"),
   679 => (x"c8",x"48",x"c0",x"86"),
   680 => (x"1e",x"73",x"87",x"cd"),
   681 => (x"1e",x"d9",x"ff",x"c0"),
   682 => (x"87",x"de",x"d7",x"ff"),
   683 => (x"d0",x"c1",x"86",x"c8"),
   684 => (x"1e",x"73",x"1e",x"d4"),
   685 => (x"c8",x"87",x"e7",x"f1"),
   686 => (x"05",x"98",x"70",x"86"),
   687 => (x"c0",x"87",x"c5",x"c0"),
   688 => (x"87",x"eb",x"c7",x"48"),
   689 => (x"1e",x"f1",x"ff",x"c0"),
   690 => (x"87",x"d0",x"d6",x"ff"),
   691 => (x"c2",x"c1",x"86",x"c4"),
   692 => (x"d6",x"ff",x"1e",x"c7"),
   693 => (x"86",x"c4",x"87",x"f4"),
   694 => (x"c2",x"c1",x"1e",x"c8"),
   695 => (x"d1",x"c1",x"1e",x"df"),
   696 => (x"ed",x"f9",x"1e",x"e6"),
   697 => (x"70",x"86",x"cc",x"87"),
   698 => (x"c9",x"c0",x"05",x"98"),
   699 => (x"dc",x"d8",x"c1",x"87"),
   700 => (x"c0",x"78",x"c1",x"48"),
   701 => (x"1e",x"c8",x"87",x"e4"),
   702 => (x"1e",x"e8",x"c2",x"c1"),
   703 => (x"1e",x"ca",x"d1",x"c1"),
   704 => (x"cc",x"87",x"cf",x"f9"),
   705 => (x"02",x"98",x"70",x"86"),
   706 => (x"c1",x"87",x"cf",x"c0"),
   707 => (x"ff",x"1e",x"d8",x"c0"),
   708 => (x"c4",x"87",x"f7",x"d5"),
   709 => (x"c6",x"48",x"c0",x"86"),
   710 => (x"d8",x"c1",x"87",x"d5"),
   711 => (x"49",x"bf",x"97",x"d2"),
   712 => (x"05",x"a9",x"d5",x"c1"),
   713 => (x"c1",x"87",x"cd",x"c0"),
   714 => (x"bf",x"97",x"d3",x"d8"),
   715 => (x"a9",x"ea",x"c2",x"49"),
   716 => (x"87",x"c5",x"c0",x"02"),
   717 => (x"f6",x"c5",x"48",x"c0"),
   718 => (x"d4",x"d0",x"c1",x"87"),
   719 => (x"c3",x"49",x"bf",x"97"),
   720 => (x"c0",x"02",x"a9",x"e9"),
   721 => (x"d0",x"c1",x"87",x"d2"),
   722 => (x"49",x"bf",x"97",x"d4"),
   723 => (x"02",x"a9",x"eb",x"c3"),
   724 => (x"c0",x"87",x"c5",x"c0"),
   725 => (x"87",x"d7",x"c5",x"48"),
   726 => (x"97",x"df",x"d0",x"c1"),
   727 => (x"99",x"71",x"49",x"bf"),
   728 => (x"87",x"cc",x"c0",x"05"),
   729 => (x"97",x"e0",x"d0",x"c1"),
   730 => (x"a9",x"c2",x"49",x"bf"),
   731 => (x"87",x"c5",x"c0",x"02"),
   732 => (x"fa",x"c4",x"48",x"c0"),
   733 => (x"e1",x"d0",x"c1",x"87"),
   734 => (x"c1",x"48",x"bf",x"97"),
   735 => (x"c1",x"58",x"d8",x"d8"),
   736 => (x"49",x"bf",x"d4",x"d8"),
   737 => (x"8a",x"c1",x"4a",x"71"),
   738 => (x"5a",x"dc",x"d8",x"c1"),
   739 => (x"1e",x"71",x"1e",x"72"),
   740 => (x"1e",x"f1",x"c2",x"c1"),
   741 => (x"87",x"f2",x"d3",x"ff"),
   742 => (x"d0",x"c1",x"86",x"cc"),
   743 => (x"49",x"bf",x"97",x"e2"),
   744 => (x"d0",x"c1",x"81",x"73"),
   745 => (x"4a",x"bf",x"97",x"e3"),
   746 => (x"48",x"72",x"32",x"c8"),
   747 => (x"d8",x"c1",x"80",x"71"),
   748 => (x"d0",x"c1",x"58",x"ec"),
   749 => (x"48",x"bf",x"97",x"e4"),
   750 => (x"58",x"c0",x"d9",x"c1"),
   751 => (x"bf",x"dc",x"d8",x"c1"),
   752 => (x"87",x"da",x"c2",x"02"),
   753 => (x"c0",x"c1",x"1e",x"c8"),
   754 => (x"d1",x"c1",x"1e",x"f5"),
   755 => (x"c1",x"f6",x"1e",x"e6"),
   756 => (x"70",x"86",x"cc",x"87"),
   757 => (x"c5",x"c0",x"02",x"98"),
   758 => (x"c3",x"48",x"c0",x"87"),
   759 => (x"d8",x"c1",x"87",x"d1"),
   760 => (x"72",x"4a",x"bf",x"d4"),
   761 => (x"c1",x"30",x"c4",x"48"),
   762 => (x"c1",x"58",x"c4",x"d9"),
   763 => (x"c1",x"5a",x"fc",x"d8"),
   764 => (x"bf",x"97",x"f9",x"d0"),
   765 => (x"c1",x"31",x"c8",x"49"),
   766 => (x"bf",x"97",x"f8",x"d0"),
   767 => (x"c1",x"81",x"73",x"4b"),
   768 => (x"bf",x"97",x"fa",x"d0"),
   769 => (x"73",x"33",x"d0",x"4b"),
   770 => (x"fb",x"d0",x"c1",x"81"),
   771 => (x"d8",x"4b",x"bf",x"97"),
   772 => (x"c1",x"81",x"73",x"33"),
   773 => (x"c1",x"59",x"c8",x"d9"),
   774 => (x"91",x"bf",x"fc",x"d8"),
   775 => (x"bf",x"e8",x"d8",x"c1"),
   776 => (x"f0",x"d8",x"c1",x"81"),
   777 => (x"c1",x"d1",x"c1",x"59"),
   778 => (x"c8",x"4b",x"bf",x"97"),
   779 => (x"c0",x"d1",x"c1",x"33"),
   780 => (x"74",x"4c",x"bf",x"97"),
   781 => (x"c2",x"d1",x"c1",x"83"),
   782 => (x"d0",x"4c",x"bf",x"97"),
   783 => (x"c1",x"83",x"74",x"34"),
   784 => (x"bf",x"97",x"c3",x"d1"),
   785 => (x"d8",x"9c",x"cf",x"4c"),
   786 => (x"c1",x"83",x"74",x"34"),
   787 => (x"c2",x"5b",x"f4",x"d8"),
   788 => (x"72",x"92",x"73",x"8b"),
   789 => (x"c1",x"80",x"71",x"48"),
   790 => (x"c1",x"58",x"f8",x"d8"),
   791 => (x"d0",x"c1",x"87",x"cf"),
   792 => (x"49",x"bf",x"97",x"e6"),
   793 => (x"d0",x"c1",x"31",x"c8"),
   794 => (x"4a",x"bf",x"97",x"e5"),
   795 => (x"d9",x"c1",x"81",x"72"),
   796 => (x"31",x"c5",x"59",x"c4"),
   797 => (x"c9",x"81",x"ff",x"c7"),
   798 => (x"fc",x"d8",x"c1",x"29"),
   799 => (x"eb",x"d0",x"c1",x"59"),
   800 => (x"c8",x"4a",x"bf",x"97"),
   801 => (x"ea",x"d0",x"c1",x"32"),
   802 => (x"73",x"4b",x"bf",x"97"),
   803 => (x"c8",x"d9",x"c1",x"82"),
   804 => (x"fc",x"d8",x"c1",x"5a"),
   805 => (x"d8",x"c1",x"92",x"bf"),
   806 => (x"c1",x"82",x"bf",x"e8"),
   807 => (x"c1",x"5a",x"f8",x"d8"),
   808 => (x"c0",x"48",x"f0",x"d8"),
   809 => (x"71",x"48",x"72",x"78"),
   810 => (x"f0",x"d8",x"c1",x"80"),
   811 => (x"f3",x"48",x"c1",x"58"),
   812 => (x"5e",x"0e",x"87",x"ea"),
   813 => (x"c1",x"0e",x"5c",x"5b"),
   814 => (x"02",x"bf",x"dc",x"d8"),
   815 => (x"cc",x"87",x"cf",x"c0"),
   816 => (x"b7",x"c7",x"4a",x"66"),
   817 => (x"4b",x"66",x"cc",x"2a"),
   818 => (x"c0",x"9b",x"ff",x"c1"),
   819 => (x"66",x"cc",x"87",x"cc"),
   820 => (x"2a",x"b7",x"c8",x"4a"),
   821 => (x"c3",x"4b",x"66",x"cc"),
   822 => (x"d0",x"c1",x"9b",x"ff"),
   823 => (x"d8",x"c1",x"1e",x"d4"),
   824 => (x"72",x"49",x"bf",x"e8"),
   825 => (x"e8",x"1e",x"71",x"81"),
   826 => (x"86",x"c8",x"87",x"f4"),
   827 => (x"c0",x"05",x"98",x"70"),
   828 => (x"48",x"c0",x"87",x"c5"),
   829 => (x"c1",x"87",x"ea",x"c0"),
   830 => (x"02",x"bf",x"dc",x"d8"),
   831 => (x"73",x"87",x"d4",x"c0"),
   832 => (x"91",x"b7",x"c4",x"49"),
   833 => (x"81",x"d4",x"d0",x"c1"),
   834 => (x"ff",x"cf",x"4c",x"69"),
   835 => (x"9c",x"ff",x"ff",x"ff"),
   836 => (x"73",x"87",x"cc",x"c0"),
   837 => (x"91",x"b7",x"c2",x"49"),
   838 => (x"81",x"d4",x"d0",x"c1"),
   839 => (x"74",x"4c",x"69",x"9f"),
   840 => (x"87",x"fa",x"f1",x"48"),
   841 => (x"5c",x"5b",x"5e",x"0e"),
   842 => (x"86",x"f4",x"0e",x"5d"),
   843 => (x"48",x"76",x"4b",x"c0"),
   844 => (x"bf",x"f0",x"d8",x"c1"),
   845 => (x"c1",x"80",x"c4",x"78"),
   846 => (x"78",x"bf",x"f4",x"d8"),
   847 => (x"bf",x"dc",x"d8",x"c1"),
   848 => (x"87",x"ca",x"c0",x"02"),
   849 => (x"bf",x"d4",x"d8",x"c1"),
   850 => (x"c0",x"31",x"c4",x"49"),
   851 => (x"d8",x"c1",x"87",x"c7"),
   852 => (x"c4",x"49",x"bf",x"f8"),
   853 => (x"59",x"a6",x"cc",x"31"),
   854 => (x"66",x"c8",x"4d",x"c0"),
   855 => (x"06",x"a8",x"c0",x"48"),
   856 => (x"75",x"87",x"f5",x"c2"),
   857 => (x"71",x"99",x"cf",x"49"),
   858 => (x"db",x"c0",x"05",x"99"),
   859 => (x"d4",x"d0",x"c1",x"87"),
   860 => (x"49",x"66",x"c8",x"1e"),
   861 => (x"cc",x"80",x"c1",x"48"),
   862 => (x"1e",x"71",x"58",x"a6"),
   863 => (x"c8",x"87",x"df",x"e6"),
   864 => (x"d4",x"d0",x"c1",x"86"),
   865 => (x"87",x"c3",x"c0",x"4b"),
   866 => (x"97",x"83",x"e0",x"c0"),
   867 => (x"99",x"71",x"49",x"6b"),
   868 => (x"87",x"fb",x"c1",x"02"),
   869 => (x"c3",x"49",x"6b",x"97"),
   870 => (x"c1",x"02",x"a9",x"e5"),
   871 => (x"49",x"73",x"87",x"f1"),
   872 => (x"69",x"97",x"81",x"cb"),
   873 => (x"71",x"99",x"d8",x"49"),
   874 => (x"e2",x"c1",x"05",x"99"),
   875 => (x"ff",x"1e",x"73",x"87"),
   876 => (x"c4",x"87",x"e9",x"ca"),
   877 => (x"c0",x"1e",x"cb",x"86"),
   878 => (x"73",x"1e",x"66",x"e4"),
   879 => (x"87",x"d2",x"ee",x"1e"),
   880 => (x"98",x"70",x"86",x"cc"),
   881 => (x"87",x"c7",x"c1",x"05"),
   882 => (x"82",x"dc",x"4a",x"73"),
   883 => (x"c4",x"49",x"66",x"dc"),
   884 => (x"73",x"79",x"6a",x"81"),
   885 => (x"dc",x"82",x"da",x"4a"),
   886 => (x"81",x"c8",x"49",x"66"),
   887 => (x"70",x"48",x"6a",x"9f"),
   888 => (x"c1",x"4c",x"71",x"79"),
   889 => (x"02",x"bf",x"dc",x"d8"),
   890 => (x"73",x"87",x"d2",x"c0"),
   891 => (x"9f",x"81",x"d4",x"49"),
   892 => (x"ff",x"c0",x"49",x"69"),
   893 => (x"4a",x"71",x"99",x"ff"),
   894 => (x"c2",x"c0",x"32",x"d0"),
   895 => (x"72",x"4a",x"c0",x"87"),
   896 => (x"70",x"80",x"6c",x"48"),
   897 => (x"48",x"66",x"dc",x"7c"),
   898 => (x"48",x"c1",x"78",x"c0"),
   899 => (x"c1",x"87",x"c0",x"c1"),
   900 => (x"ad",x"66",x"c8",x"85"),
   901 => (x"87",x"cb",x"fd",x"04"),
   902 => (x"bf",x"dc",x"d8",x"c1"),
   903 => (x"87",x"ed",x"c0",x"02"),
   904 => (x"cd",x"fa",x"1e",x"6e"),
   905 => (x"c4",x"86",x"c4",x"87"),
   906 => (x"49",x"6e",x"58",x"a6"),
   907 => (x"ff",x"ff",x"ff",x"cf"),
   908 => (x"02",x"a9",x"99",x"f8"),
   909 => (x"6e",x"87",x"d6",x"c0"),
   910 => (x"c1",x"89",x"c2",x"49"),
   911 => (x"91",x"bf",x"d4",x"d8"),
   912 => (x"bf",x"ec",x"d8",x"c1"),
   913 => (x"c8",x"80",x"71",x"48"),
   914 => (x"cb",x"fc",x"58",x"a6"),
   915 => (x"f4",x"48",x"c0",x"87"),
   916 => (x"87",x"c8",x"ed",x"8e"),
   917 => (x"0e",x"5b",x"5e",x"0e"),
   918 => (x"49",x"bf",x"66",x"c8"),
   919 => (x"66",x"c8",x"81",x"c1"),
   920 => (x"c1",x"09",x"79",x"09"),
   921 => (x"99",x"bf",x"d8",x"d8"),
   922 => (x"c0",x"05",x"99",x"71"),
   923 => (x"66",x"c8",x"87",x"d0"),
   924 => (x"6b",x"83",x"c8",x"4b"),
   925 => (x"87",x"fa",x"f8",x"1e"),
   926 => (x"49",x"70",x"86",x"c4"),
   927 => (x"48",x"c1",x"7b",x"71"),
   928 => (x"0e",x"87",x"dd",x"ec"),
   929 => (x"d8",x"c1",x"0e",x"5e"),
   930 => (x"c4",x"49",x"bf",x"ec"),
   931 => (x"82",x"c8",x"4a",x"66"),
   932 => (x"8a",x"c2",x"4a",x"6a"),
   933 => (x"bf",x"d4",x"d8",x"c1"),
   934 => (x"c1",x"81",x"72",x"92"),
   935 => (x"4a",x"bf",x"d8",x"d8"),
   936 => (x"9a",x"bf",x"66",x"c4"),
   937 => (x"66",x"c8",x"81",x"72"),
   938 => (x"e1",x"1e",x"71",x"1e"),
   939 => (x"86",x"c8",x"87",x"f0"),
   940 => (x"c0",x"05",x"98",x"70"),
   941 => (x"48",x"c0",x"87",x"c5"),
   942 => (x"c1",x"87",x"c2",x"c0"),
   943 => (x"87",x"e2",x"eb",x"48"),
   944 => (x"5c",x"5b",x"5e",x"0e"),
   945 => (x"1e",x"66",x"cc",x"0e"),
   946 => (x"1e",x"cc",x"d9",x"c1"),
   947 => (x"c8",x"87",x"d5",x"f9"),
   948 => (x"02",x"98",x"70",x"86"),
   949 => (x"c1",x"87",x"d4",x"c1"),
   950 => (x"49",x"bf",x"d0",x"d9"),
   951 => (x"c9",x"81",x"ff",x"c7"),
   952 => (x"c0",x"4c",x"71",x"29"),
   953 => (x"c2",x"fd",x"c0",x"4b"),
   954 => (x"ef",x"c5",x"ff",x"1e"),
   955 => (x"c0",x"86",x"c4",x"87"),
   956 => (x"c1",x"06",x"ac",x"b7"),
   957 => (x"66",x"d0",x"87",x"c7"),
   958 => (x"cc",x"d9",x"c1",x"1e"),
   959 => (x"87",x"c3",x"fe",x"1e"),
   960 => (x"98",x"70",x"86",x"c8"),
   961 => (x"87",x"c5",x"c0",x"05"),
   962 => (x"f2",x"c0",x"48",x"c0"),
   963 => (x"cc",x"d9",x"c1",x"87"),
   964 => (x"87",x"c0",x"fd",x"1e"),
   965 => (x"66",x"d0",x"86",x"c4"),
   966 => (x"80",x"c0",x"c8",x"48"),
   967 => (x"c1",x"58",x"a6",x"d4"),
   968 => (x"ab",x"b7",x"74",x"83"),
   969 => (x"87",x"ce",x"ff",x"04"),
   970 => (x"cc",x"87",x"d2",x"c0"),
   971 => (x"fd",x"c0",x"1e",x"66"),
   972 => (x"c5",x"ff",x"1e",x"db"),
   973 => (x"86",x"c8",x"87",x"d4"),
   974 => (x"c2",x"c0",x"48",x"c0"),
   975 => (x"e9",x"48",x"c1",x"87"),
   976 => (x"70",x"4f",x"87",x"dc"),
   977 => (x"64",x"65",x"6e",x"65"),
   978 => (x"6c",x"69",x"66",x"20"),
   979 => (x"6c",x"20",x"2c",x"65"),
   980 => (x"69",x"64",x"61",x"6f"),
   981 => (x"2e",x"2e",x"67",x"6e"),
   982 => (x"43",x"00",x"0a",x"2e"),
   983 => (x"74",x"27",x"6e",x"61"),
   984 => (x"65",x"70",x"6f",x"20"),
   985 => (x"73",x"25",x"20",x"6e"),
   986 => (x"65",x"52",x"00",x"0a"),
   987 => (x"6f",x"20",x"64",x"61"),
   988 => (x"42",x"4d",x"20",x"66"),
   989 => (x"61",x"66",x"20",x"52"),
   990 => (x"64",x"65",x"6c",x"69"),
   991 => (x"6f",x"4e",x"00",x"0a"),
   992 => (x"72",x"61",x"70",x"20"),
   993 => (x"69",x"74",x"69",x"74"),
   994 => (x"73",x"20",x"6e",x"6f"),
   995 => (x"61",x"6e",x"67",x"69"),
   996 => (x"65",x"72",x"75",x"74"),
   997 => (x"75",x"6f",x"66",x"20"),
   998 => (x"00",x"0a",x"64",x"6e"),
   999 => (x"73",x"52",x"42",x"4d"),
  1000 => (x"3a",x"65",x"7a",x"69"),
  1001 => (x"2c",x"64",x"25",x"20"),
  1002 => (x"72",x"61",x"70",x"20"),
  1003 => (x"69",x"74",x"69",x"74"),
  1004 => (x"69",x"73",x"6e",x"6f"),
  1005 => (x"20",x"3a",x"65",x"7a"),
  1006 => (x"20",x"2c",x"64",x"25"),
  1007 => (x"73",x"66",x"66",x"6f"),
  1008 => (x"6f",x"20",x"74",x"65"),
  1009 => (x"69",x"73",x"20",x"66"),
  1010 => (x"25",x"20",x"3a",x"67"),
  1011 => (x"73",x"20",x"2c",x"64"),
  1012 => (x"30",x"20",x"67",x"69"),
  1013 => (x"0a",x"78",x"25",x"78"),
  1014 => (x"61",x"65",x"52",x"00"),
  1015 => (x"67",x"6e",x"69",x"64"),
  1016 => (x"6f",x"6f",x"62",x"20"),
  1017 => (x"65",x"73",x"20",x"74"),
  1018 => (x"72",x"6f",x"74",x"63"),
  1019 => (x"0a",x"64",x"25",x"20"),
  1020 => (x"61",x"65",x"52",x"00"),
  1021 => (x"6f",x"62",x"20",x"64"),
  1022 => (x"73",x"20",x"74",x"6f"),
  1023 => (x"6f",x"74",x"63",x"65"),
  1024 => (x"72",x"66",x"20",x"72"),
  1025 => (x"66",x"20",x"6d",x"6f"),
  1026 => (x"74",x"73",x"72",x"69"),
  1027 => (x"72",x"61",x"70",x"20"),
  1028 => (x"69",x"74",x"69",x"74"),
  1029 => (x"00",x"0a",x"6e",x"6f"),
  1030 => (x"75",x"73",x"6e",x"55"),
  1031 => (x"72",x"6f",x"70",x"70"),
  1032 => (x"20",x"64",x"65",x"74"),
  1033 => (x"74",x"72",x"61",x"70"),
  1034 => (x"6f",x"69",x"74",x"69"),
  1035 => (x"79",x"74",x"20",x"6e"),
  1036 => (x"0d",x"21",x"65",x"70"),
  1037 => (x"54",x"41",x"46",x"00"),
  1038 => (x"20",x"20",x"32",x"33"),
  1039 => (x"65",x"52",x"00",x"20"),
  1040 => (x"6e",x"69",x"64",x"61"),
  1041 => (x"42",x"4d",x"20",x"67"),
  1042 => (x"4d",x"00",x"0a",x"52"),
  1043 => (x"73",x"20",x"52",x"42"),
  1044 => (x"65",x"63",x"63",x"75"),
  1045 => (x"75",x"66",x"73",x"73"),
  1046 => (x"20",x"79",x"6c",x"6c"),
  1047 => (x"64",x"61",x"65",x"72"),
  1048 => (x"41",x"46",x"00",x"0a"),
  1049 => (x"20",x"36",x"31",x"54"),
  1050 => (x"46",x"00",x"20",x"20"),
  1051 => (x"32",x"33",x"54",x"41"),
  1052 => (x"00",x"20",x"20",x"20"),
  1053 => (x"74",x"72",x"61",x"50"),
  1054 => (x"6f",x"69",x"74",x"69"),
  1055 => (x"75",x"6f",x"63",x"6e"),
  1056 => (x"25",x"20",x"74",x"6e"),
  1057 => (x"48",x"00",x"0a",x"64"),
  1058 => (x"69",x"74",x"6e",x"75"),
  1059 => (x"66",x"20",x"67",x"6e"),
  1060 => (x"66",x"20",x"72",x"6f"),
  1061 => (x"73",x"65",x"6c",x"69"),
  1062 => (x"65",x"74",x"73",x"79"),
  1063 => (x"46",x"00",x"0a",x"6d"),
  1064 => (x"32",x"33",x"54",x"41"),
  1065 => (x"00",x"20",x"20",x"20"),
  1066 => (x"31",x"54",x"41",x"46"),
  1067 => (x"20",x"20",x"20",x"36"),
  1068 => (x"75",x"6c",x"43",x"00"),
  1069 => (x"72",x"65",x"74",x"73"),
  1070 => (x"7a",x"69",x"73",x"20"),
  1071 => (x"25",x"20",x"3a",x"65"),
  1072 => (x"43",x"20",x"2c",x"64"),
  1073 => (x"74",x"73",x"75",x"6c"),
  1074 => (x"6d",x"20",x"72",x"65"),
  1075 => (x"2c",x"6b",x"73",x"61"),
  1076 => (x"0a",x"64",x"25",x"20"),
  1077 => (x"0e",x"5e",x"0e",x"00"),
  1078 => (x"d8",x"49",x"66",x"c4"),
  1079 => (x"99",x"ff",x"c3",x"29"),
  1080 => (x"c8",x"4a",x"66",x"c4"),
  1081 => (x"c0",x"fc",x"cf",x"2a"),
  1082 => (x"c4",x"b1",x"72",x"9a"),
  1083 => (x"32",x"c8",x"4a",x"66"),
  1084 => (x"c0",x"f0",x"ff",x"c0"),
  1085 => (x"b1",x"72",x"9a",x"c0"),
  1086 => (x"d8",x"4a",x"66",x"c4"),
  1087 => (x"c0",x"c0",x"ff",x"32"),
  1088 => (x"72",x"9a",x"c0",x"c0"),
  1089 => (x"c6",x"48",x"71",x"b1"),
  1090 => (x"26",x"4d",x"26",x"87"),
  1091 => (x"26",x"4b",x"26",x"4c"),
  1092 => (x"0e",x"5e",x"0e",x"4f"),
  1093 => (x"c8",x"4a",x"66",x"c4"),
  1094 => (x"9a",x"ff",x"c3",x"2a"),
  1095 => (x"9a",x"ff",x"ff",x"cf"),
  1096 => (x"c8",x"49",x"66",x"c4"),
  1097 => (x"c0",x"fc",x"cf",x"31"),
  1098 => (x"cf",x"b1",x"72",x"99"),
  1099 => (x"71",x"99",x"ff",x"ff"),
  1100 => (x"87",x"db",x"ff",x"48"),
  1101 => (x"c4",x"0e",x"5e",x"0e"),
  1102 => (x"29",x"d0",x"49",x"66"),
  1103 => (x"99",x"ff",x"ff",x"cf"),
  1104 => (x"d0",x"4a",x"66",x"c4"),
  1105 => (x"c0",x"c0",x"f0",x"32"),
  1106 => (x"71",x"b1",x"72",x"9a"),
  1107 => (x"87",x"ff",x"fe",x"48"),
  1108 => (x"c8",x"0e",x"5e",x"0e"),
  1109 => (x"49",x"72",x"4a",x"66"),
  1110 => (x"99",x"71",x"8a",x"c1"),
  1111 => (x"c4",x"87",x"de",x"02"),
  1112 => (x"48",x"bf",x"97",x"66"),
  1113 => (x"b8",x"80",x"c0",x"fe"),
  1114 => (x"08",x"78",x"08",x"fc"),
  1115 => (x"c1",x"48",x"66",x"c4"),
  1116 => (x"58",x"a6",x"c8",x"80"),
  1117 => (x"8a",x"c1",x"49",x"72"),
  1118 => (x"e2",x"05",x"99",x"71"),
  1119 => (x"26",x"87",x"c6",x"87"),
  1120 => (x"26",x"4c",x"26",x"4d"),
  1121 => (x"0e",x"4f",x"26",x"4b"),
  1122 => (x"c8",x"0e",x"5b",x"5e"),
  1123 => (x"d9",x"c1",x"1e",x"66"),
  1124 => (x"cf",x"ee",x"1e",x"cc"),
  1125 => (x"70",x"86",x"c8",x"87"),
  1126 => (x"e1",x"c1",x"02",x"98"),
  1127 => (x"d0",x"d9",x"c1",x"87"),
  1128 => (x"cf",x"c1",x"4b",x"bf"),
  1129 => (x"fa",x"fe",x"1e",x"c8"),
  1130 => (x"86",x"c4",x"87",x"f2"),
  1131 => (x"78",x"c1",x"48",x"f8"),
  1132 => (x"c1",x"02",x"9b",x"73"),
  1133 => (x"d0",x"c1",x"87",x"c2"),
  1134 => (x"d9",x"c1",x"1e",x"d4"),
  1135 => (x"c2",x"f3",x"1e",x"cc"),
  1136 => (x"70",x"86",x"c8",x"87"),
  1137 => (x"87",x"c5",x"05",x"98"),
  1138 => (x"c4",x"c1",x"48",x"c0"),
  1139 => (x"cc",x"d9",x"c1",x"87"),
  1140 => (x"87",x"c0",x"f2",x"1e"),
  1141 => (x"c0",x"c8",x"86",x"c4"),
  1142 => (x"c6",x"04",x"ab",x"b7"),
  1143 => (x"49",x"c0",x"c8",x"87"),
  1144 => (x"73",x"87",x"c4",x"8b"),
  1145 => (x"71",x"4b",x"c0",x"49"),
  1146 => (x"d4",x"d0",x"c1",x"1e"),
  1147 => (x"87",x"e0",x"fd",x"1e"),
  1148 => (x"9b",x"73",x"86",x"c8"),
  1149 => (x"87",x"fe",x"fe",x"05"),
  1150 => (x"78",x"c0",x"48",x"f8"),
  1151 => (x"66",x"c8",x"87",x"d1"),
  1152 => (x"e1",x"cf",x"c1",x"1e"),
  1153 => (x"c1",x"fa",x"fe",x"1e"),
  1154 => (x"c0",x"86",x"c8",x"87"),
  1155 => (x"c1",x"87",x"c2",x"48"),
  1156 => (x"87",x"ef",x"fd",x"48"),
  1157 => (x"c1",x"49",x"c0",x"1e"),
  1158 => (x"b7",x"c0",x"d0",x"81"),
  1159 => (x"f6",x"ff",x"04",x"a9"),
  1160 => (x"87",x"e1",x"fd",x"87"),
  1161 => (x"5c",x"5b",x"5e",x"0e"),
  1162 => (x"ff",x"1e",x"0e",x"5d"),
  1163 => (x"ce",x"c1",x"4d",x"d4"),
  1164 => (x"f8",x"fe",x"1e",x"cc"),
  1165 => (x"86",x"c4",x"87",x"e6"),
  1166 => (x"48",x"e4",x"d9",x"c1"),
  1167 => (x"d0",x"ff",x"50",x"c0"),
  1168 => (x"c0",x"c8",x"48",x"bf"),
  1169 => (x"a6",x"c4",x"98",x"c0"),
  1170 => (x"d0",x"02",x"6e",x"58"),
  1171 => (x"bf",x"d0",x"ff",x"87"),
  1172 => (x"c0",x"c0",x"c8",x"48"),
  1173 => (x"58",x"a6",x"c4",x"98"),
  1174 => (x"f0",x"ff",x"05",x"6e"),
  1175 => (x"48",x"d0",x"ff",x"87"),
  1176 => (x"d4",x"78",x"e1",x"c0"),
  1177 => (x"c3",x"4b",x"c0",x"7d"),
  1178 => (x"4c",x"6d",x"7d",x"ff"),
  1179 => (x"c1",x"02",x"9c",x"74"),
  1180 => (x"d9",x"c1",x"87",x"f7"),
  1181 => (x"81",x"73",x"49",x"e4"),
  1182 => (x"ff",x"c3",x"51",x"74"),
  1183 => (x"87",x"d4",x"fe",x"98"),
  1184 => (x"f6",x"fe",x"1e",x"74"),
  1185 => (x"86",x"c4",x"87",x"f6"),
  1186 => (x"05",x"ac",x"fb",x"c0"),
  1187 => (x"c8",x"87",x"cd",x"c1"),
  1188 => (x"d4",x"03",x"ab",x"b7"),
  1189 => (x"e4",x"d9",x"c1",x"87"),
  1190 => (x"c0",x"81",x"73",x"49"),
  1191 => (x"83",x"c1",x"51",x"e0"),
  1192 => (x"04",x"ab",x"b7",x"c8"),
  1193 => (x"d5",x"87",x"ee",x"ff"),
  1194 => (x"ab",x"b7",x"c8",x"87"),
  1195 => (x"87",x"ce",x"c0",x"06"),
  1196 => (x"48",x"ea",x"d9",x"c1"),
  1197 => (x"c1",x"50",x"fe",x"c1"),
  1198 => (x"c0",x"48",x"eb",x"d9"),
  1199 => (x"d9",x"c1",x"50",x"f1"),
  1200 => (x"d2",x"c1",x"48",x"ec"),
  1201 => (x"ed",x"d9",x"c1",x"50"),
  1202 => (x"50",x"cf",x"c1",x"48"),
  1203 => (x"48",x"ee",x"d9",x"c1"),
  1204 => (x"c1",x"50",x"cd",x"c1"),
  1205 => (x"c0",x"48",x"ef",x"d9"),
  1206 => (x"87",x"cd",x"c0",x"50"),
  1207 => (x"ff",x"c3",x"83",x"c1"),
  1208 => (x"74",x"4c",x"6d",x"7d"),
  1209 => (x"c9",x"fe",x"05",x"9c"),
  1210 => (x"7d",x"ff",x"c3",x"87"),
  1211 => (x"cb",x"c0",x"02",x"6d"),
  1212 => (x"7d",x"ff",x"c3",x"87"),
  1213 => (x"99",x"71",x"49",x"6d"),
  1214 => (x"87",x"f5",x"ff",x"05"),
  1215 => (x"48",x"bf",x"d0",x"ff"),
  1216 => (x"98",x"c0",x"c0",x"c8"),
  1217 => (x"6e",x"58",x"a6",x"c4"),
  1218 => (x"87",x"d0",x"c0",x"02"),
  1219 => (x"48",x"bf",x"d0",x"ff"),
  1220 => (x"98",x"c0",x"c0",x"c8"),
  1221 => (x"6e",x"58",x"a6",x"c4"),
  1222 => (x"87",x"f0",x"ff",x"05"),
  1223 => (x"c0",x"48",x"d0",x"ff"),
  1224 => (x"ef",x"fb",x"78",x"e0"),
  1225 => (x"e4",x"d9",x"c1",x"87"),
  1226 => (x"ef",x"f4",x"fe",x"1e"),
  1227 => (x"c1",x"86",x"c4",x"87"),
  1228 => (x"fe",x"1e",x"e2",x"ce"),
  1229 => (x"c4",x"87",x"e5",x"f4"),
  1230 => (x"e6",x"c5",x"ff",x"86"),
  1231 => (x"02",x"98",x"70",x"87"),
  1232 => (x"ff",x"87",x"cf",x"c0"),
  1233 => (x"70",x"87",x"dd",x"d9"),
  1234 => (x"c5",x"c0",x"02",x"98"),
  1235 => (x"c0",x"49",x"c1",x"87"),
  1236 => (x"49",x"c0",x"87",x"c2"),
  1237 => (x"c0",x"02",x"99",x"71"),
  1238 => (x"d9",x"c1",x"87",x"dc"),
  1239 => (x"e6",x"f8",x"1e",x"e4"),
  1240 => (x"70",x"86",x"c4",x"87"),
  1241 => (x"cd",x"c0",x"02",x"98"),
  1242 => (x"c6",x"ce",x"c1",x"87"),
  1243 => (x"eb",x"f3",x"fe",x"1e"),
  1244 => (x"c0",x"86",x"c4",x"87"),
  1245 => (x"ce",x"c1",x"87",x"ca"),
  1246 => (x"f3",x"fe",x"1e",x"f8"),
  1247 => (x"86",x"c4",x"87",x"de"),
  1248 => (x"f7",x"26",x"48",x"c0"),
  1249 => (x"6f",x"44",x"87",x"f9"),
  1250 => (x"00",x"0a",x"65",x"6e"),
  1251 => (x"63",x"74",x"65",x"46"),
  1252 => (x"67",x"6e",x"69",x"68"),
  1253 => (x"6e",x"6f",x"63",x"20"),
  1254 => (x"74",x"73",x"20",x"66"),
  1255 => (x"67",x"6e",x"69",x"72"),
  1256 => (x"6e",x"49",x"00",x"0a"),
  1257 => (x"61",x"69",x"74",x"69"),
  1258 => (x"69",x"7a",x"69",x"6c"),
  1259 => (x"53",x"20",x"67",x"6e"),
  1260 => (x"61",x"63",x"20",x"44"),
  1261 => (x"00",x"0a",x"64",x"72"),
  1262 => (x"62",x"20",x"44",x"53"),
  1263 => (x"20",x"74",x"6f",x"6f"),
  1264 => (x"6c",x"69",x"61",x"66"),
  1265 => (x"00",x"0a",x"64",x"65"),
  1266 => (x"6e",x"65",x"70",x"4f"),
  1267 => (x"66",x"20",x"64",x"65"),
  1268 => (x"2c",x"65",x"6c",x"69"),
  1269 => (x"61",x"6f",x"6c",x"20"),
  1270 => (x"67",x"6e",x"69",x"64"),
  1271 => (x"0a",x"2e",x"2e",x"2e"),
  1272 => (x"6e",x"61",x"43",x"00"),
  1273 => (x"6f",x"20",x"74",x"27"),
  1274 => (x"20",x"6e",x"65",x"70"),
  1275 => (x"00",x"0a",x"73",x"25"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
