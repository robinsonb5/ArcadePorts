
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Boot_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of Boot_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f8",x"eb",x"c1",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"f8",x"eb",x"c1"),
    18 => (x"48",x"cc",x"e2",x"c1"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"c9",x"e2",x"c1",x"87"),
    25 => (x"c5",x"e2",x"c1",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"d0",x"c1",x"87",x"f7"),
    29 => (x"e2",x"c1",x"87",x"f4"),
    30 => (x"e2",x"c1",x"4d",x"c9"),
    31 => (x"ad",x"74",x"4c",x"c9"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"fc",x"98",x"00",x"87"),
    35 => (x"5b",x"5e",x"0e",x"87"),
    36 => (x"f8",x"0e",x"5d",x"5c"),
    37 => (x"c0",x"4c",x"71",x"86"),
    38 => (x"c1",x"4d",x"66",x"e4"),
    39 => (x"4b",x"a7",x"ed",x"df"),
    40 => (x"7e",x"a7",x"cd",x"c2"),
    41 => (x"c0",x"48",x"a6",x"c4"),
    42 => (x"05",x"9c",x"74",x"78"),
    43 => (x"f0",x"c0",x"87",x"c6"),
    44 => (x"87",x"c6",x"c1",x"53"),
    45 => (x"c0",x"02",x"9c",x"74"),
    46 => (x"49",x"74",x"87",x"e2"),
    47 => (x"4a",x"66",x"dc",x"1e"),
    48 => (x"71",x"87",x"c9",x"cb"),
    49 => (x"6e",x"49",x"26",x"4a"),
    50 => (x"d8",x"53",x"12",x"82"),
    51 => (x"fb",x"ca",x"4a",x"66"),
    52 => (x"4c",x"49",x"70",x"87"),
    53 => (x"9c",x"74",x"8d",x"c1"),
    54 => (x"87",x"de",x"ff",x"05"),
    55 => (x"06",x"ad",x"b7",x"c0"),
    56 => (x"e8",x"c0",x"87",x"d8"),
    57 => (x"87",x"c5",x"02",x"66"),
    58 => (x"c3",x"4a",x"f0",x"c0"),
    59 => (x"4a",x"e0",x"c0",x"87"),
    60 => (x"8d",x"c1",x"53",x"72"),
    61 => (x"01",x"ad",x"b7",x"c0"),
    62 => (x"de",x"c1",x"87",x"e8"),
    63 => (x"02",x"ab",x"a7",x"ce"),
    64 => (x"dc",x"87",x"e0",x"c0"),
    65 => (x"e0",x"c0",x"4c",x"66"),
    66 => (x"8b",x"c1",x"1e",x"66"),
    67 => (x"74",x"49",x"6b",x"97"),
    68 => (x"66",x"86",x"c4",x"0f"),
    69 => (x"c8",x"80",x"c1",x"48"),
    70 => (x"dd",x"c1",x"58",x"a6"),
    71 => (x"05",x"ab",x"a7",x"ee"),
    72 => (x"c4",x"87",x"e3",x"ff"),
    73 => (x"8e",x"f8",x"48",x"66"),
    74 => (x"4c",x"26",x"4d",x"26"),
    75 => (x"4f",x"26",x"4b",x"26"),
    76 => (x"33",x"32",x"31",x"30"),
    77 => (x"37",x"36",x"35",x"34"),
    78 => (x"42",x"41",x"39",x"38"),
    79 => (x"46",x"45",x"44",x"43"),
    80 => (x"5b",x"5e",x"0e",x"00"),
    81 => (x"71",x"0e",x"5d",x"5c"),
    82 => (x"13",x"4d",x"ff",x"4b"),
    83 => (x"d7",x"02",x"9c",x"4c"),
    84 => (x"d4",x"85",x"c1",x"87"),
    85 => (x"49",x"74",x"1e",x"66"),
    86 => (x"c4",x"0f",x"66",x"d4"),
    87 => (x"05",x"a8",x"74",x"86"),
    88 => (x"4c",x"13",x"87",x"c6"),
    89 => (x"87",x"e9",x"05",x"9c"),
    90 => (x"4d",x"26",x"48",x"75"),
    91 => (x"4b",x"26",x"4c",x"26"),
    92 => (x"5e",x"0e",x"4f",x"26"),
    93 => (x"0e",x"5d",x"5c",x"5b"),
    94 => (x"a6",x"c8",x"86",x"e8"),
    95 => (x"66",x"e8",x"c0",x"59"),
    96 => (x"c8",x"4c",x"c0",x"4d"),
    97 => (x"78",x"c0",x"48",x"a6"),
    98 => (x"bf",x"97",x"66",x"c4"),
    99 => (x"48",x"66",x"c4",x"4b"),
   100 => (x"a6",x"c8",x"80",x"c1"),
   101 => (x"02",x"9b",x"73",x"58"),
   102 => (x"c8",x"87",x"d3",x"c6"),
   103 => (x"d9",x"c5",x"02",x"66"),
   104 => (x"48",x"a6",x"cc",x"87"),
   105 => (x"80",x"fc",x"78",x"c0"),
   106 => (x"4a",x"73",x"78",x"c0"),
   107 => (x"02",x"8a",x"e0",x"c0"),
   108 => (x"c3",x"87",x"c8",x"c3"),
   109 => (x"c2",x"c3",x"02",x"8a"),
   110 => (x"02",x"8a",x"c2",x"87"),
   111 => (x"8a",x"87",x"ea",x"c2"),
   112 => (x"87",x"f7",x"c2",x"02"),
   113 => (x"c2",x"02",x"8a",x"c4"),
   114 => (x"8a",x"c2",x"87",x"f1"),
   115 => (x"87",x"eb",x"c2",x"02"),
   116 => (x"c2",x"02",x"8a",x"c3"),
   117 => (x"8a",x"d4",x"87",x"ed"),
   118 => (x"87",x"fa",x"c0",x"02"),
   119 => (x"c5",x"c1",x"02",x"8a"),
   120 => (x"02",x"8a",x"ca",x"87"),
   121 => (x"c1",x"87",x"f7",x"c0"),
   122 => (x"e5",x"c1",x"02",x"8a"),
   123 => (x"c0",x"02",x"8a",x"87"),
   124 => (x"8a",x"c5",x"87",x"e4"),
   125 => (x"c3",x"87",x"df",x"02"),
   126 => (x"cd",x"c1",x"02",x"8a"),
   127 => (x"02",x"8a",x"c4",x"87"),
   128 => (x"c3",x"87",x"e3",x"c0"),
   129 => (x"e5",x"c0",x"02",x"8a"),
   130 => (x"02",x"8a",x"c2",x"87"),
   131 => (x"8a",x"c3",x"87",x"c8"),
   132 => (x"c1",x"87",x"d3",x"02"),
   133 => (x"a6",x"cc",x"87",x"f9"),
   134 => (x"c2",x"78",x"ca",x"48"),
   135 => (x"a6",x"cc",x"87",x"d2"),
   136 => (x"c2",x"78",x"c2",x"48"),
   137 => (x"a6",x"cc",x"87",x"ca"),
   138 => (x"c2",x"78",x"d0",x"48"),
   139 => (x"f0",x"c0",x"87",x"c2"),
   140 => (x"f0",x"c0",x"1e",x"66"),
   141 => (x"85",x"c4",x"1e",x"66"),
   142 => (x"8a",x"c4",x"4a",x"75"),
   143 => (x"c0",x"fc",x"49",x"6a"),
   144 => (x"70",x"86",x"c8",x"87"),
   145 => (x"c1",x"4c",x"a4",x"49"),
   146 => (x"a6",x"c8",x"87",x"e6"),
   147 => (x"c1",x"78",x"c1",x"48"),
   148 => (x"f0",x"c0",x"87",x"de"),
   149 => (x"85",x"c4",x"1e",x"66"),
   150 => (x"8a",x"c4",x"4a",x"75"),
   151 => (x"f0",x"c0",x"49",x"6a"),
   152 => (x"86",x"c4",x"0f",x"66"),
   153 => (x"c7",x"c1",x"84",x"c1"),
   154 => (x"66",x"f0",x"c0",x"87"),
   155 => (x"49",x"e5",x"c0",x"1e"),
   156 => (x"0f",x"66",x"f0",x"c0"),
   157 => (x"84",x"c1",x"86",x"c4"),
   158 => (x"c8",x"87",x"f5",x"c0"),
   159 => (x"78",x"c1",x"48",x"a6"),
   160 => (x"d0",x"87",x"ed",x"c0"),
   161 => (x"78",x"c1",x"48",x"a6"),
   162 => (x"78",x"c1",x"80",x"f8"),
   163 => (x"c0",x"87",x"e1",x"c0"),
   164 => (x"db",x"06",x"ab",x"f0"),
   165 => (x"ab",x"f9",x"c0",x"87"),
   166 => (x"d4",x"87",x"d5",x"03"),
   167 => (x"92",x"ca",x"4a",x"66"),
   168 => (x"f0",x"c0",x"49",x"73"),
   169 => (x"49",x"a1",x"72",x"89"),
   170 => (x"48",x"59",x"a6",x"d8"),
   171 => (x"78",x"c1",x"80",x"f4"),
   172 => (x"c1",x"02",x"66",x"cc"),
   173 => (x"85",x"c4",x"87",x"e5"),
   174 => (x"89",x"c4",x"49",x"75"),
   175 => (x"e4",x"c1",x"7e",x"69"),
   176 => (x"87",x"d5",x"05",x"ab"),
   177 => (x"b7",x"c0",x"48",x"6e"),
   178 => (x"87",x"cd",x"03",x"a8"),
   179 => (x"c1",x"49",x"ed",x"c0"),
   180 => (x"48",x"6e",x"87",x"fb"),
   181 => (x"70",x"88",x"08",x"c0"),
   182 => (x"1e",x"66",x"d0",x"7e"),
   183 => (x"c0",x"1e",x"66",x"d8"),
   184 => (x"c0",x"1e",x"66",x"f8"),
   185 => (x"dc",x"1e",x"66",x"f8"),
   186 => (x"d4",x"1e",x"49",x"66"),
   187 => (x"dc",x"f6",x"49",x"66"),
   188 => (x"70",x"86",x"d4",x"87"),
   189 => (x"c0",x"4c",x"a4",x"49"),
   190 => (x"e5",x"c0",x"87",x"e1"),
   191 => (x"87",x"cf",x"05",x"ab"),
   192 => (x"c0",x"48",x"a6",x"d0"),
   193 => (x"c0",x"80",x"c4",x"78"),
   194 => (x"c1",x"80",x"f4",x"78"),
   195 => (x"c0",x"87",x"cc",x"78"),
   196 => (x"73",x"1e",x"66",x"f0"),
   197 => (x"66",x"f0",x"c0",x"49"),
   198 => (x"c4",x"86",x"c4",x"0f"),
   199 => (x"4b",x"bf",x"97",x"66"),
   200 => (x"c1",x"48",x"66",x"c4"),
   201 => (x"58",x"a6",x"c8",x"80"),
   202 => (x"f9",x"05",x"9b",x"73"),
   203 => (x"48",x"74",x"87",x"ed"),
   204 => (x"4d",x"26",x"8e",x"e8"),
   205 => (x"4b",x"26",x"4c",x"26"),
   206 => (x"c0",x"1e",x"4f",x"26"),
   207 => (x"1e",x"a7",x"ce",x"1e"),
   208 => (x"d0",x"1e",x"a6",x"d0"),
   209 => (x"e9",x"f8",x"49",x"66"),
   210 => (x"26",x"8e",x"f4",x"87"),
   211 => (x"86",x"fc",x"1e",x"4f"),
   212 => (x"c0",x"ff",x"4a",x"71"),
   213 => (x"c4",x"48",x"69",x"49"),
   214 => (x"7e",x"70",x"98",x"c0"),
   215 => (x"f4",x"02",x"98",x"48"),
   216 => (x"48",x"79",x"72",x"87"),
   217 => (x"4f",x"26",x"8e",x"fc"),
   218 => (x"5c",x"5b",x"5e",x"0e"),
   219 => (x"c0",x"4b",x"71",x"0e"),
   220 => (x"9a",x"4a",x"13",x"4c"),
   221 => (x"72",x"87",x"cd",x"02"),
   222 => (x"87",x"d1",x"ff",x"49"),
   223 => (x"4a",x"13",x"84",x"c1"),
   224 => (x"87",x"f3",x"05",x"9a"),
   225 => (x"4c",x"26",x"48",x"74"),
   226 => (x"4f",x"26",x"4b",x"26"),
   227 => (x"72",x"1e",x"73",x"1e"),
   228 => (x"e7",x"c0",x"02",x"9a"),
   229 => (x"c1",x"48",x"c0",x"87"),
   230 => (x"06",x"a9",x"72",x"4b"),
   231 => (x"82",x"72",x"87",x"d1"),
   232 => (x"73",x"87",x"c9",x"06"),
   233 => (x"01",x"a9",x"72",x"83"),
   234 => (x"87",x"c3",x"87",x"f4"),
   235 => (x"72",x"3a",x"b2",x"c1"),
   236 => (x"73",x"89",x"03",x"a9"),
   237 => (x"2a",x"c1",x"07",x"80"),
   238 => (x"87",x"f3",x"05",x"2b"),
   239 => (x"4f",x"26",x"4b",x"26"),
   240 => (x"c4",x"1e",x"75",x"1e"),
   241 => (x"a1",x"b7",x"71",x"4d"),
   242 => (x"c1",x"b9",x"ff",x"04"),
   243 => (x"07",x"bd",x"c3",x"81"),
   244 => (x"04",x"a2",x"b7",x"72"),
   245 => (x"82",x"c1",x"ba",x"ff"),
   246 => (x"fe",x"07",x"bd",x"c1"),
   247 => (x"2d",x"c1",x"87",x"ee"),
   248 => (x"c1",x"b8",x"ff",x"04"),
   249 => (x"04",x"2d",x"07",x"80"),
   250 => (x"81",x"c1",x"b9",x"ff"),
   251 => (x"26",x"4d",x"26",x"07"),
   252 => (x"dc",x"ff",x"1e",x"4f"),
   253 => (x"4a",x"d4",x"ff",x"86"),
   254 => (x"6a",x"7a",x"ff",x"c3"),
   255 => (x"7a",x"ff",x"c3",x"49"),
   256 => (x"30",x"c8",x"48",x"6a"),
   257 => (x"a6",x"c8",x"7e",x"70"),
   258 => (x"48",x"66",x"c4",x"59"),
   259 => (x"a6",x"cc",x"b0",x"6e"),
   260 => (x"c3",x"49",x"70",x"58"),
   261 => (x"48",x"6a",x"7a",x"ff"),
   262 => (x"58",x"a6",x"30",x"d0"),
   263 => (x"d0",x"59",x"a6",x"d4"),
   264 => (x"66",x"cc",x"48",x"66"),
   265 => (x"58",x"a6",x"d8",x"b0"),
   266 => (x"ff",x"c3",x"49",x"70"),
   267 => (x"d8",x"48",x"6a",x"7a"),
   268 => (x"58",x"a6",x"dc",x"30"),
   269 => (x"59",x"a6",x"e0",x"c0"),
   270 => (x"d8",x"48",x"66",x"dc"),
   271 => (x"e4",x"c0",x"b0",x"66"),
   272 => (x"ff",x"70",x"58",x"a6"),
   273 => (x"4f",x"26",x"8e",x"dc"),
   274 => (x"ff",x"86",x"e8",x"1e"),
   275 => (x"ff",x"c3",x"4a",x"d4"),
   276 => (x"c3",x"49",x"6a",x"7a"),
   277 => (x"31",x"c8",x"7a",x"ff"),
   278 => (x"48",x"6a",x"7e",x"71"),
   279 => (x"a6",x"c8",x"b0",x"6e"),
   280 => (x"c3",x"49",x"70",x"58"),
   281 => (x"31",x"c8",x"7a",x"ff"),
   282 => (x"6a",x"59",x"a6",x"cc"),
   283 => (x"b0",x"66",x"c8",x"48"),
   284 => (x"70",x"58",x"a6",x"d0"),
   285 => (x"7a",x"ff",x"c3",x"49"),
   286 => (x"a6",x"d4",x"31",x"c8"),
   287 => (x"d0",x"48",x"6a",x"59"),
   288 => (x"a6",x"d8",x"b0",x"66"),
   289 => (x"8e",x"e8",x"70",x"58"),
   290 => (x"5e",x"0e",x"4f",x"26"),
   291 => (x"0e",x"5d",x"5c",x"5b"),
   292 => (x"d4",x"ff",x"4a",x"71"),
   293 => (x"c3",x"49",x"72",x"4d"),
   294 => (x"7d",x"71",x"99",x"ff"),
   295 => (x"bf",x"e0",x"e2",x"c1"),
   296 => (x"d0",x"87",x"c8",x"05"),
   297 => (x"30",x"c9",x"48",x"66"),
   298 => (x"d0",x"58",x"a6",x"d4"),
   299 => (x"29",x"d8",x"49",x"66"),
   300 => (x"71",x"99",x"ff",x"c3"),
   301 => (x"49",x"66",x"d0",x"7d"),
   302 => (x"ff",x"c3",x"29",x"d0"),
   303 => (x"d0",x"7d",x"71",x"99"),
   304 => (x"29",x"c8",x"49",x"66"),
   305 => (x"71",x"99",x"ff",x"c3"),
   306 => (x"49",x"66",x"d0",x"7d"),
   307 => (x"71",x"99",x"ff",x"c3"),
   308 => (x"d0",x"49",x"72",x"7d"),
   309 => (x"99",x"ff",x"c3",x"29"),
   310 => (x"4b",x"6d",x"7d",x"71"),
   311 => (x"4c",x"ff",x"f0",x"c9"),
   312 => (x"05",x"ab",x"ff",x"c3"),
   313 => (x"ff",x"c3",x"87",x"d0"),
   314 => (x"c1",x"4b",x"6d",x"7d"),
   315 => (x"87",x"c6",x"02",x"8c"),
   316 => (x"02",x"ab",x"ff",x"c3"),
   317 => (x"48",x"73",x"87",x"f0"),
   318 => (x"4c",x"26",x"4d",x"26"),
   319 => (x"4f",x"26",x"4b",x"26"),
   320 => (x"ff",x"49",x"c0",x"1e"),
   321 => (x"ff",x"c3",x"48",x"d4"),
   322 => (x"c3",x"81",x"c1",x"78"),
   323 => (x"04",x"a9",x"b7",x"c8"),
   324 => (x"4f",x"26",x"87",x"f1"),
   325 => (x"e7",x"1e",x"73",x"1e"),
   326 => (x"df",x"f8",x"c4",x"87"),
   327 => (x"c0",x"1e",x"c0",x"4b"),
   328 => (x"f7",x"c1",x"f0",x"ff"),
   329 => (x"87",x"e2",x"fd",x"49"),
   330 => (x"a8",x"c1",x"86",x"c4"),
   331 => (x"87",x"ea",x"c0",x"05"),
   332 => (x"c3",x"48",x"d4",x"ff"),
   333 => (x"c0",x"c1",x"78",x"ff"),
   334 => (x"c0",x"c0",x"c0",x"c0"),
   335 => (x"f0",x"e1",x"c0",x"1e"),
   336 => (x"fd",x"49",x"e9",x"c1"),
   337 => (x"86",x"c4",x"87",x"c4"),
   338 => (x"ca",x"05",x"98",x"70"),
   339 => (x"48",x"d4",x"ff",x"87"),
   340 => (x"c1",x"78",x"ff",x"c3"),
   341 => (x"fe",x"87",x"cb",x"48"),
   342 => (x"8b",x"c1",x"87",x"e6"),
   343 => (x"87",x"fd",x"fe",x"05"),
   344 => (x"d7",x"fe",x"48",x"c0"),
   345 => (x"1e",x"73",x"1e",x"87"),
   346 => (x"c3",x"48",x"d4",x"ff"),
   347 => (x"e0",x"d6",x"78",x"ff"),
   348 => (x"87",x"f4",x"f7",x"49"),
   349 => (x"1e",x"c0",x"4b",x"d3"),
   350 => (x"c1",x"f0",x"ff",x"c0"),
   351 => (x"c9",x"fc",x"49",x"c1"),
   352 => (x"70",x"86",x"c4",x"87"),
   353 => (x"87",x"ca",x"05",x"98"),
   354 => (x"c3",x"48",x"d4",x"ff"),
   355 => (x"48",x"c1",x"78",x"ff"),
   356 => (x"eb",x"fd",x"87",x"cb"),
   357 => (x"05",x"8b",x"c1",x"87"),
   358 => (x"c0",x"87",x"db",x"ff"),
   359 => (x"87",x"dc",x"fd",x"48"),
   360 => (x"00",x"44",x"4d",x"43"),
   361 => (x"5c",x"5b",x"5e",x"0e"),
   362 => (x"d4",x"ff",x"0e",x"5d"),
   363 => (x"87",x"d0",x"fd",x"4d"),
   364 => (x"c0",x"1e",x"ea",x"c6"),
   365 => (x"c8",x"c1",x"f0",x"e1"),
   366 => (x"87",x"ce",x"fb",x"49"),
   367 => (x"da",x"1e",x"4b",x"70"),
   368 => (x"f5",x"f5",x"1e",x"e3"),
   369 => (x"c1",x"86",x"cc",x"87"),
   370 => (x"87",x"c8",x"02",x"ab"),
   371 => (x"c0",x"87",x"d6",x"fe"),
   372 => (x"87",x"ca",x"c2",x"48"),
   373 => (x"70",x"87",x"f1",x"f9"),
   374 => (x"ff",x"ff",x"cf",x"49"),
   375 => (x"a9",x"ea",x"c6",x"99"),
   376 => (x"fd",x"87",x"c8",x"02"),
   377 => (x"48",x"c0",x"87",x"ff"),
   378 => (x"c3",x"87",x"f3",x"c1"),
   379 => (x"f1",x"c0",x"7d",x"ff"),
   380 => (x"87",x"e0",x"fc",x"4c"),
   381 => (x"c1",x"02",x"98",x"70"),
   382 => (x"1e",x"c0",x"87",x"cb"),
   383 => (x"c1",x"f0",x"ff",x"c0"),
   384 => (x"c5",x"fa",x"49",x"fa"),
   385 => (x"70",x"86",x"c4",x"87"),
   386 => (x"c0",x"05",x"9b",x"4b"),
   387 => (x"d9",x"1e",x"87",x"ed"),
   388 => (x"e5",x"f4",x"1e",x"e1"),
   389 => (x"7d",x"ff",x"c3",x"87"),
   390 => (x"d9",x"1e",x"4b",x"6d"),
   391 => (x"d9",x"f4",x"1e",x"ed"),
   392 => (x"c3",x"86",x"d0",x"87"),
   393 => (x"7d",x"7d",x"7d",x"ff"),
   394 => (x"c1",x"49",x"73",x"7d"),
   395 => (x"c5",x"02",x"99",x"c0"),
   396 => (x"c0",x"48",x"c1",x"87"),
   397 => (x"48",x"c0",x"87",x"e8"),
   398 => (x"73",x"87",x"e3",x"c0"),
   399 => (x"1e",x"fb",x"d9",x"1e"),
   400 => (x"c8",x"87",x"f7",x"f3"),
   401 => (x"05",x"ac",x"c2",x"86"),
   402 => (x"c7",x"da",x"87",x"cc"),
   403 => (x"87",x"ea",x"f3",x"1e"),
   404 => (x"48",x"c0",x"86",x"c4"),
   405 => (x"8c",x"c1",x"87",x"c8"),
   406 => (x"87",x"d5",x"fe",x"05"),
   407 => (x"d7",x"fa",x"48",x"c0"),
   408 => (x"44",x"4d",x"43",x"87"),
   409 => (x"25",x"20",x"38",x"35"),
   410 => (x"20",x"20",x"0a",x"64"),
   411 => (x"44",x"4d",x"43",x"00"),
   412 => (x"32",x"5f",x"38",x"35"),
   413 => (x"0a",x"64",x"25",x"20"),
   414 => (x"43",x"00",x"20",x"20"),
   415 => (x"38",x"35",x"44",x"4d"),
   416 => (x"0a",x"64",x"25",x"20"),
   417 => (x"53",x"00",x"20",x"20"),
   418 => (x"20",x"43",x"48",x"44"),
   419 => (x"74",x"69",x"6e",x"49"),
   420 => (x"69",x"6c",x"61",x"69"),
   421 => (x"69",x"74",x"61",x"7a"),
   422 => (x"65",x"20",x"6e",x"6f"),
   423 => (x"72",x"6f",x"72",x"72"),
   424 => (x"63",x"00",x"0a",x"21"),
   425 => (x"43",x"5f",x"64",x"6d"),
   426 => (x"20",x"38",x"44",x"4d"),
   427 => (x"70",x"73",x"65",x"72"),
   428 => (x"65",x"73",x"6e",x"6f"),
   429 => (x"64",x"25",x"20",x"3a"),
   430 => (x"5e",x"0e",x"00",x"0a"),
   431 => (x"0e",x"5d",x"5c",x"5b"),
   432 => (x"4d",x"d0",x"ff",x"1e"),
   433 => (x"4b",x"c0",x"c0",x"c8"),
   434 => (x"48",x"e0",x"e2",x"c1"),
   435 => (x"cb",x"de",x"78",x"c1"),
   436 => (x"87",x"d4",x"f2",x"49"),
   437 => (x"48",x"6d",x"4c",x"c7"),
   438 => (x"7e",x"70",x"98",x"73"),
   439 => (x"cb",x"02",x"98",x"48"),
   440 => (x"73",x"48",x"6d",x"87"),
   441 => (x"48",x"7e",x"70",x"98"),
   442 => (x"87",x"f5",x"05",x"98"),
   443 => (x"cf",x"f8",x"7d",x"c2"),
   444 => (x"73",x"48",x"6d",x"87"),
   445 => (x"48",x"7e",x"70",x"98"),
   446 => (x"87",x"cb",x"02",x"98"),
   447 => (x"98",x"73",x"48",x"6d"),
   448 => (x"98",x"48",x"7e",x"70"),
   449 => (x"c3",x"87",x"f5",x"05"),
   450 => (x"c0",x"1e",x"c0",x"7d"),
   451 => (x"c0",x"c1",x"d0",x"e5"),
   452 => (x"87",x"f6",x"f5",x"49"),
   453 => (x"a8",x"c1",x"86",x"c4"),
   454 => (x"4c",x"87",x"c1",x"05"),
   455 => (x"cb",x"05",x"ac",x"c2"),
   456 => (x"49",x"c6",x"de",x"87"),
   457 => (x"c0",x"87",x"c1",x"f1"),
   458 => (x"87",x"d6",x"c1",x"48"),
   459 => (x"fe",x"05",x"8c",x"c1"),
   460 => (x"ef",x"f9",x"87",x"e4"),
   461 => (x"e4",x"e2",x"c1",x"87"),
   462 => (x"05",x"98",x"70",x"58"),
   463 => (x"1e",x"c1",x"87",x"cd"),
   464 => (x"c1",x"f0",x"ff",x"c0"),
   465 => (x"c1",x"f5",x"49",x"d0"),
   466 => (x"ff",x"86",x"c4",x"87"),
   467 => (x"ff",x"c3",x"48",x"d4"),
   468 => (x"87",x"fa",x"c5",x"78"),
   469 => (x"58",x"e8",x"e2",x"c1"),
   470 => (x"cf",x"de",x"1e",x"70"),
   471 => (x"87",x"da",x"ef",x"1e"),
   472 => (x"48",x"6d",x"86",x"c8"),
   473 => (x"7e",x"70",x"98",x"73"),
   474 => (x"cb",x"02",x"98",x"48"),
   475 => (x"73",x"48",x"6d",x"87"),
   476 => (x"48",x"7e",x"70",x"98"),
   477 => (x"87",x"f5",x"05",x"98"),
   478 => (x"d4",x"ff",x"7d",x"c2"),
   479 => (x"78",x"ff",x"c3",x"48"),
   480 => (x"f5",x"26",x"48",x"c1"),
   481 => (x"45",x"49",x"87",x"f2"),
   482 => (x"53",x"00",x"52",x"52"),
   483 => (x"53",x"00",x"49",x"50"),
   484 => (x"61",x"63",x"20",x"44"),
   485 => (x"73",x"20",x"64",x"72"),
   486 => (x"20",x"65",x"7a",x"69"),
   487 => (x"25",x"20",x"73",x"69"),
   488 => (x"0e",x"00",x"0a",x"64"),
   489 => (x"5d",x"5c",x"5b",x"5e"),
   490 => (x"d0",x"4b",x"71",x"0e"),
   491 => (x"4c",x"c0",x"4d",x"66"),
   492 => (x"df",x"cd",x"ee",x"c5"),
   493 => (x"48",x"d4",x"ff",x"4a"),
   494 => (x"68",x"78",x"ff",x"c3"),
   495 => (x"a9",x"fe",x"c3",x"49"),
   496 => (x"87",x"ca",x"c1",x"05"),
   497 => (x"48",x"dc",x"e2",x"c1"),
   498 => (x"b7",x"c4",x"78",x"c0"),
   499 => (x"87",x"d8",x"04",x"ad"),
   500 => (x"70",x"87",x"de",x"f0"),
   501 => (x"e2",x"c1",x"43",x"49"),
   502 => (x"71",x"48",x"bf",x"dc"),
   503 => (x"e0",x"e2",x"c1",x"80"),
   504 => (x"b7",x"8d",x"c4",x"58"),
   505 => (x"87",x"e8",x"03",x"ad"),
   506 => (x"06",x"ad",x"b7",x"c0"),
   507 => (x"d4",x"ff",x"87",x"dd"),
   508 => (x"78",x"ff",x"c3",x"48"),
   509 => (x"c1",x"53",x"49",x"68"),
   510 => (x"48",x"bf",x"dc",x"e2"),
   511 => (x"e2",x"c1",x"80",x"71"),
   512 => (x"8d",x"c1",x"58",x"e0"),
   513 => (x"01",x"ad",x"b7",x"c0"),
   514 => (x"c1",x"87",x"e3",x"ff"),
   515 => (x"8a",x"c1",x"4c",x"4a"),
   516 => (x"87",x"e1",x"fe",x"05"),
   517 => (x"c3",x"48",x"d4",x"ff"),
   518 => (x"48",x"74",x"78",x"ff"),
   519 => (x"0e",x"87",x"d9",x"f3"),
   520 => (x"5d",x"5c",x"5b",x"5e"),
   521 => (x"4b",x"71",x"1e",x"0e"),
   522 => (x"4d",x"c0",x"c0",x"c8"),
   523 => (x"d4",x"ff",x"4c",x"c0"),
   524 => (x"78",x"ff",x"c3",x"48"),
   525 => (x"48",x"bf",x"d0",x"ff"),
   526 => (x"7e",x"70",x"98",x"75"),
   527 => (x"cd",x"02",x"98",x"48"),
   528 => (x"bf",x"d0",x"ff",x"87"),
   529 => (x"70",x"98",x"75",x"48"),
   530 => (x"05",x"98",x"48",x"7e"),
   531 => (x"d0",x"ff",x"87",x"f3"),
   532 => (x"78",x"c3",x"c4",x"48"),
   533 => (x"c3",x"48",x"d4",x"ff"),
   534 => (x"1e",x"73",x"78",x"ff"),
   535 => (x"c1",x"f0",x"ff",x"c0"),
   536 => (x"e5",x"f0",x"49",x"d1"),
   537 => (x"70",x"86",x"c4",x"87"),
   538 => (x"cf",x"02",x"9a",x"4a"),
   539 => (x"1e",x"73",x"1e",x"87"),
   540 => (x"1e",x"ee",x"e2",x"c0"),
   541 => (x"cc",x"87",x"c3",x"eb"),
   542 => (x"87",x"ec",x"c0",x"86"),
   543 => (x"d8",x"1e",x"c0",x"c8"),
   544 => (x"de",x"fc",x"49",x"66"),
   545 => (x"70",x"86",x"c4",x"87"),
   546 => (x"bf",x"d0",x"ff",x"4c"),
   547 => (x"70",x"98",x"75",x"48"),
   548 => (x"02",x"98",x"48",x"7e"),
   549 => (x"d0",x"ff",x"87",x"cd"),
   550 => (x"98",x"75",x"48",x"bf"),
   551 => (x"98",x"48",x"7e",x"70"),
   552 => (x"ff",x"87",x"f3",x"05"),
   553 => (x"78",x"c2",x"48",x"d0"),
   554 => (x"f1",x"26",x"48",x"74"),
   555 => (x"65",x"52",x"87",x"ca"),
   556 => (x"63",x"20",x"64",x"61"),
   557 => (x"61",x"6d",x"6d",x"6f"),
   558 => (x"66",x"20",x"64",x"6e"),
   559 => (x"65",x"6c",x"69",x"61"),
   560 => (x"74",x"61",x"20",x"64"),
   561 => (x"20",x"64",x"25",x"20"),
   562 => (x"29",x"64",x"25",x"28"),
   563 => (x"5e",x"0e",x"00",x"0a"),
   564 => (x"0e",x"5d",x"5c",x"5b"),
   565 => (x"c0",x"1e",x"c0",x"1e"),
   566 => (x"c9",x"c1",x"f0",x"ff"),
   567 => (x"87",x"ea",x"ee",x"49"),
   568 => (x"e2",x"c1",x"1e",x"d2"),
   569 => (x"fa",x"fa",x"49",x"e8"),
   570 => (x"c0",x"86",x"c8",x"87"),
   571 => (x"d2",x"85",x"c1",x"4d"),
   572 => (x"f8",x"04",x"ad",x"b7"),
   573 => (x"e8",x"e2",x"c1",x"87"),
   574 => (x"c3",x"49",x"bf",x"97"),
   575 => (x"c0",x"c1",x"99",x"c0"),
   576 => (x"e7",x"c0",x"05",x"a9"),
   577 => (x"ef",x"e2",x"c1",x"87"),
   578 => (x"d0",x"49",x"bf",x"97"),
   579 => (x"f0",x"e2",x"c1",x"31"),
   580 => (x"c8",x"4a",x"bf",x"97"),
   581 => (x"c1",x"b1",x"72",x"32"),
   582 => (x"bf",x"97",x"f1",x"e2"),
   583 => (x"4d",x"71",x"b1",x"4a"),
   584 => (x"ff",x"ff",x"ff",x"cf"),
   585 => (x"ca",x"85",x"c1",x"9d"),
   586 => (x"87",x"e3",x"c2",x"35"),
   587 => (x"97",x"f1",x"e2",x"c1"),
   588 => (x"33",x"c1",x"4b",x"bf"),
   589 => (x"e2",x"c1",x"9b",x"c6"),
   590 => (x"49",x"bf",x"97",x"f2"),
   591 => (x"71",x"29",x"b7",x"c7"),
   592 => (x"ed",x"e2",x"c1",x"b3"),
   593 => (x"48",x"49",x"bf",x"97"),
   594 => (x"7e",x"70",x"98",x"cf"),
   595 => (x"97",x"ee",x"e2",x"c1"),
   596 => (x"9c",x"c3",x"4c",x"bf"),
   597 => (x"e2",x"c1",x"34",x"ca"),
   598 => (x"49",x"bf",x"97",x"ef"),
   599 => (x"b4",x"71",x"31",x"c2"),
   600 => (x"97",x"f0",x"e2",x"c1"),
   601 => (x"c0",x"c3",x"49",x"bf"),
   602 => (x"29",x"b7",x"c6",x"99"),
   603 => (x"1e",x"74",x"b4",x"71"),
   604 => (x"73",x"1e",x"66",x"c4"),
   605 => (x"d5",x"e7",x"c0",x"1e"),
   606 => (x"87",x"fe",x"e6",x"1e"),
   607 => (x"48",x"c1",x"83",x"c2"),
   608 => (x"4b",x"70",x"30",x"73"),
   609 => (x"c2",x"e8",x"c0",x"1e"),
   610 => (x"87",x"ee",x"e6",x"1e"),
   611 => (x"66",x"d8",x"48",x"c1"),
   612 => (x"58",x"a6",x"dc",x"30"),
   613 => (x"4d",x"49",x"a4",x"c1"),
   614 => (x"66",x"d8",x"95",x"73"),
   615 => (x"c0",x"1e",x"75",x"1e"),
   616 => (x"e6",x"1e",x"cb",x"e8"),
   617 => (x"e4",x"c0",x"87",x"d4"),
   618 => (x"c8",x"48",x"6e",x"86"),
   619 => (x"06",x"a8",x"b7",x"c0"),
   620 => (x"35",x"c1",x"87",x"d2"),
   621 => (x"b7",x"c1",x"48",x"6e"),
   622 => (x"48",x"7e",x"70",x"28"),
   623 => (x"a8",x"b7",x"c0",x"c8"),
   624 => (x"87",x"ee",x"ff",x"01"),
   625 => (x"e8",x"c0",x"1e",x"75"),
   626 => (x"ed",x"e5",x"1e",x"e1"),
   627 => (x"75",x"86",x"c8",x"87"),
   628 => (x"e3",x"ec",x"26",x"48"),
   629 => (x"73",x"5f",x"63",x"87"),
   630 => (x"5f",x"65",x"7a",x"69"),
   631 => (x"74",x"6c",x"75",x"6d"),
   632 => (x"64",x"25",x"20",x"3a"),
   633 => (x"65",x"72",x"20",x"2c"),
   634 => (x"62",x"5f",x"64",x"61"),
   635 => (x"65",x"6c",x"5f",x"6c"),
   636 => (x"25",x"20",x"3a",x"6e"),
   637 => (x"63",x"20",x"2c",x"64"),
   638 => (x"65",x"7a",x"69",x"73"),
   639 => (x"64",x"25",x"20",x"3a"),
   640 => (x"75",x"4d",x"00",x"0a"),
   641 => (x"25",x"20",x"74",x"6c"),
   642 => (x"25",x"00",x"0a",x"64"),
   643 => (x"6c",x"62",x"20",x"64"),
   644 => (x"73",x"6b",x"63",x"6f"),
   645 => (x"20",x"66",x"6f",x"20"),
   646 => (x"65",x"7a",x"69",x"73"),
   647 => (x"0a",x"64",x"25",x"20"),
   648 => (x"20",x"64",x"25",x"00"),
   649 => (x"63",x"6f",x"6c",x"62"),
   650 => (x"6f",x"20",x"73",x"6b"),
   651 => (x"31",x"35",x"20",x"66"),
   652 => (x"79",x"62",x"20",x"32"),
   653 => (x"0a",x"73",x"65",x"74"),
   654 => (x"5b",x"5e",x"0e",x"00"),
   655 => (x"4b",x"71",x"0e",x"5c"),
   656 => (x"66",x"d0",x"4c",x"c0"),
   657 => (x"a8",x"b7",x"c0",x"48"),
   658 => (x"87",x"eb",x"c0",x"06"),
   659 => (x"c0",x"fe",x"4a",x"13"),
   660 => (x"66",x"cc",x"ba",x"82"),
   661 => (x"fe",x"49",x"bf",x"97"),
   662 => (x"cc",x"b9",x"81",x"c0"),
   663 => (x"80",x"c1",x"48",x"66"),
   664 => (x"71",x"58",x"a6",x"d0"),
   665 => (x"c4",x"02",x"aa",x"b7"),
   666 => (x"cc",x"48",x"c1",x"87"),
   667 => (x"d0",x"84",x"c1",x"87"),
   668 => (x"04",x"ac",x"b7",x"66"),
   669 => (x"c0",x"87",x"d5",x"ff"),
   670 => (x"26",x"87",x"c2",x"48"),
   671 => (x"26",x"4c",x"26",x"4d"),
   672 => (x"0e",x"4f",x"26",x"4b"),
   673 => (x"5d",x"5c",x"5b",x"5e"),
   674 => (x"c2",x"eb",x"c1",x"0e"),
   675 => (x"c0",x"78",x"c0",x"48"),
   676 => (x"e3",x"49",x"dc",x"f9"),
   677 => (x"e2",x"c1",x"87",x"d2"),
   678 => (x"49",x"c0",x"1e",x"fa"),
   679 => (x"c4",x"87",x"c0",x"f6"),
   680 => (x"05",x"98",x"70",x"86"),
   681 => (x"f6",x"c0",x"87",x"cc"),
   682 => (x"fb",x"e2",x"49",x"c8"),
   683 => (x"cb",x"48",x"c0",x"87"),
   684 => (x"f9",x"c0",x"87",x"d3"),
   685 => (x"ef",x"e2",x"49",x"e9"),
   686 => (x"c1",x"4b",x"c0",x"87"),
   687 => (x"c1",x"48",x"e6",x"eb"),
   688 => (x"c0",x"1e",x"c8",x"78"),
   689 => (x"c1",x"1e",x"c0",x"fa"),
   690 => (x"fd",x"49",x"f0",x"e3"),
   691 => (x"86",x"c8",x"87",x"eb"),
   692 => (x"c6",x"05",x"98",x"70"),
   693 => (x"e6",x"eb",x"c1",x"87"),
   694 => (x"c8",x"78",x"c0",x"48"),
   695 => (x"c9",x"fa",x"c0",x"1e"),
   696 => (x"cc",x"e4",x"c1",x"1e"),
   697 => (x"87",x"d1",x"fd",x"49"),
   698 => (x"98",x"70",x"86",x"c8"),
   699 => (x"c1",x"87",x"c6",x"05"),
   700 => (x"c0",x"48",x"e6",x"eb"),
   701 => (x"e6",x"eb",x"c1",x"78"),
   702 => (x"fa",x"c0",x"1e",x"bf"),
   703 => (x"f9",x"e0",x"1e",x"d2"),
   704 => (x"c1",x"86",x"c8",x"87"),
   705 => (x"02",x"bf",x"e6",x"eb"),
   706 => (x"c1",x"87",x"cc",x"c2"),
   707 => (x"48",x"4d",x"fa",x"e2"),
   708 => (x"4c",x"a0",x"fe",x"c6"),
   709 => (x"9f",x"f8",x"ea",x"c1"),
   710 => (x"c7",x"1e",x"49",x"bf"),
   711 => (x"48",x"49",x"a0",x"fe"),
   712 => (x"89",x"a0",x"c2",x"f8"),
   713 => (x"1e",x"d0",x"1e",x"71"),
   714 => (x"c0",x"1e",x"c0",x"c8"),
   715 => (x"e0",x"1e",x"fa",x"f6"),
   716 => (x"86",x"d4",x"87",x"c8"),
   717 => (x"69",x"49",x"a4",x"c8"),
   718 => (x"f8",x"ea",x"c1",x"4b"),
   719 => (x"c5",x"49",x"bf",x"9f"),
   720 => (x"05",x"a9",x"ea",x"d6"),
   721 => (x"c8",x"87",x"cc",x"c0"),
   722 => (x"49",x"6a",x"4a",x"a4"),
   723 => (x"70",x"87",x"c9",x"d6"),
   724 => (x"c7",x"87",x"dc",x"4b"),
   725 => (x"9f",x"49",x"a5",x"fe"),
   726 => (x"e9",x"ca",x"49",x"69"),
   727 => (x"c0",x"02",x"a9",x"d5"),
   728 => (x"f6",x"c0",x"87",x"cd"),
   729 => (x"df",x"ff",x"49",x"dc"),
   730 => (x"48",x"c0",x"87",x"fe"),
   731 => (x"73",x"87",x"d6",x"c8"),
   732 => (x"f7",x"f7",x"c0",x"1e"),
   733 => (x"c1",x"df",x"ff",x"1e"),
   734 => (x"fa",x"e2",x"c1",x"87"),
   735 => (x"f2",x"49",x"73",x"1e"),
   736 => (x"86",x"cc",x"87",x"dd"),
   737 => (x"c0",x"05",x"98",x"70"),
   738 => (x"48",x"c0",x"87",x"c5"),
   739 => (x"c0",x"87",x"f6",x"c7"),
   740 => (x"ff",x"49",x"cf",x"f8"),
   741 => (x"c0",x"87",x"d1",x"df"),
   742 => (x"ff",x"1e",x"e5",x"fa"),
   743 => (x"c8",x"87",x"db",x"de"),
   744 => (x"fd",x"fa",x"c0",x"1e"),
   745 => (x"cc",x"e4",x"c1",x"1e"),
   746 => (x"87",x"cd",x"fa",x"49"),
   747 => (x"98",x"70",x"86",x"cc"),
   748 => (x"87",x"c9",x"c0",x"05"),
   749 => (x"48",x"c2",x"eb",x"c1"),
   750 => (x"e4",x"c0",x"78",x"c1"),
   751 => (x"c0",x"1e",x"c8",x"87"),
   752 => (x"c1",x"1e",x"c6",x"fb"),
   753 => (x"f9",x"49",x"f0",x"e3"),
   754 => (x"86",x"c8",x"87",x"ef"),
   755 => (x"c0",x"02",x"98",x"70"),
   756 => (x"f8",x"c0",x"87",x"cf"),
   757 => (x"dd",x"ff",x"1e",x"f6"),
   758 => (x"86",x"c4",x"87",x"e0"),
   759 => (x"e4",x"c6",x"48",x"c0"),
   760 => (x"f8",x"ea",x"c1",x"87"),
   761 => (x"c1",x"49",x"bf",x"97"),
   762 => (x"c0",x"05",x"a9",x"d5"),
   763 => (x"ea",x"c1",x"87",x"cd"),
   764 => (x"49",x"bf",x"97",x"f9"),
   765 => (x"02",x"a9",x"ea",x"c2"),
   766 => (x"c0",x"87",x"c5",x"c0"),
   767 => (x"87",x"c5",x"c6",x"48"),
   768 => (x"97",x"fa",x"e2",x"c1"),
   769 => (x"e9",x"c3",x"49",x"bf"),
   770 => (x"d2",x"c0",x"02",x"a9"),
   771 => (x"fa",x"e2",x"c1",x"87"),
   772 => (x"c3",x"49",x"bf",x"97"),
   773 => (x"c0",x"02",x"a9",x"eb"),
   774 => (x"48",x"c0",x"87",x"c5"),
   775 => (x"c1",x"87",x"e6",x"c5"),
   776 => (x"bf",x"97",x"c5",x"e3"),
   777 => (x"c0",x"05",x"99",x"49"),
   778 => (x"e3",x"c1",x"87",x"cc"),
   779 => (x"49",x"bf",x"97",x"c6"),
   780 => (x"c0",x"02",x"a9",x"c2"),
   781 => (x"48",x"c0",x"87",x"c5"),
   782 => (x"c1",x"87",x"ca",x"c5"),
   783 => (x"bf",x"97",x"c7",x"e3"),
   784 => (x"fe",x"ea",x"c1",x"48"),
   785 => (x"4a",x"49",x"70",x"58"),
   786 => (x"eb",x"c1",x"8a",x"c1"),
   787 => (x"1e",x"72",x"5a",x"c2"),
   788 => (x"fb",x"c0",x"1e",x"71"),
   789 => (x"db",x"ff",x"1e",x"cf"),
   790 => (x"86",x"cc",x"87",x"e0"),
   791 => (x"97",x"c8",x"e3",x"c1"),
   792 => (x"81",x"73",x"49",x"bf"),
   793 => (x"97",x"c9",x"e3",x"c1"),
   794 => (x"32",x"c8",x"4a",x"bf"),
   795 => (x"48",x"c6",x"eb",x"c1"),
   796 => (x"c1",x"78",x"a1",x"72"),
   797 => (x"bf",x"97",x"ca",x"e3"),
   798 => (x"de",x"eb",x"c1",x"48"),
   799 => (x"c2",x"eb",x"c1",x"58"),
   800 => (x"e6",x"c2",x"02",x"bf"),
   801 => (x"c0",x"1e",x"c8",x"87"),
   802 => (x"c1",x"1e",x"d3",x"f9"),
   803 => (x"f6",x"49",x"cc",x"e4"),
   804 => (x"86",x"c8",x"87",x"e7"),
   805 => (x"c0",x"02",x"98",x"70"),
   806 => (x"48",x"c0",x"87",x"c5"),
   807 => (x"c1",x"87",x"e6",x"c3"),
   808 => (x"4a",x"bf",x"fa",x"ea"),
   809 => (x"c1",x"30",x"c4",x"48"),
   810 => (x"c1",x"58",x"e2",x"eb"),
   811 => (x"c1",x"5a",x"da",x"eb"),
   812 => (x"bf",x"97",x"df",x"e3"),
   813 => (x"c1",x"31",x"c8",x"49"),
   814 => (x"bf",x"97",x"de",x"e3"),
   815 => (x"c1",x"49",x"a1",x"4b"),
   816 => (x"bf",x"97",x"e0",x"e3"),
   817 => (x"73",x"33",x"d0",x"4b"),
   818 => (x"e3",x"c1",x"49",x"a1"),
   819 => (x"4b",x"bf",x"97",x"e1"),
   820 => (x"a1",x"73",x"33",x"d8"),
   821 => (x"e6",x"eb",x"c1",x"49"),
   822 => (x"e2",x"eb",x"c1",x"59"),
   823 => (x"eb",x"c1",x"49",x"bf"),
   824 => (x"c1",x"91",x"bf",x"da"),
   825 => (x"81",x"bf",x"c6",x"eb"),
   826 => (x"59",x"ce",x"eb",x"c1"),
   827 => (x"97",x"e7",x"e3",x"c1"),
   828 => (x"33",x"c8",x"4b",x"bf"),
   829 => (x"97",x"e6",x"e3",x"c1"),
   830 => (x"4b",x"a3",x"4c",x"bf"),
   831 => (x"97",x"e8",x"e3",x"c1"),
   832 => (x"34",x"d0",x"4c",x"bf"),
   833 => (x"c1",x"4b",x"a3",x"74"),
   834 => (x"bf",x"97",x"e9",x"e3"),
   835 => (x"d8",x"9c",x"cf",x"4c"),
   836 => (x"4b",x"a3",x"74",x"34"),
   837 => (x"5b",x"d2",x"eb",x"c1"),
   838 => (x"bf",x"ce",x"eb",x"c1"),
   839 => (x"73",x"8b",x"c2",x"4b"),
   840 => (x"d2",x"eb",x"c1",x"92"),
   841 => (x"78",x"a1",x"72",x"48"),
   842 => (x"c1",x"87",x"d8",x"c1"),
   843 => (x"bf",x"97",x"cc",x"e3"),
   844 => (x"c1",x"31",x"c8",x"49"),
   845 => (x"bf",x"97",x"cb",x"e3"),
   846 => (x"c1",x"49",x"a1",x"4a"),
   847 => (x"c1",x"59",x"e2",x"eb"),
   848 => (x"49",x"bf",x"de",x"eb"),
   849 => (x"ff",x"c7",x"31",x"c5"),
   850 => (x"c1",x"29",x"c9",x"81"),
   851 => (x"c1",x"59",x"da",x"eb"),
   852 => (x"bf",x"97",x"d1",x"e3"),
   853 => (x"c1",x"32",x"c8",x"4a"),
   854 => (x"bf",x"97",x"d0",x"e3"),
   855 => (x"c1",x"4a",x"a2",x"4b"),
   856 => (x"c1",x"5a",x"e6",x"eb"),
   857 => (x"4a",x"bf",x"e2",x"eb"),
   858 => (x"bf",x"da",x"eb",x"c1"),
   859 => (x"c6",x"eb",x"c1",x"92"),
   860 => (x"eb",x"c1",x"82",x"bf"),
   861 => (x"eb",x"c1",x"5a",x"d6"),
   862 => (x"78",x"c0",x"48",x"ce"),
   863 => (x"48",x"ca",x"eb",x"c1"),
   864 => (x"c1",x"78",x"a1",x"72"),
   865 => (x"87",x"f3",x"f3",x"48"),
   866 => (x"64",x"61",x"65",x"52"),
   867 => (x"20",x"66",x"6f",x"20"),
   868 => (x"20",x"52",x"42",x"4d"),
   869 => (x"6c",x"69",x"61",x"66"),
   870 => (x"00",x"0a",x"64",x"65"),
   871 => (x"70",x"20",x"6f",x"4e"),
   872 => (x"69",x"74",x"72",x"61"),
   873 => (x"6e",x"6f",x"69",x"74"),
   874 => (x"67",x"69",x"73",x"20"),
   875 => (x"75",x"74",x"61",x"6e"),
   876 => (x"66",x"20",x"65",x"72"),
   877 => (x"64",x"6e",x"75",x"6f"),
   878 => (x"42",x"4d",x"00",x"0a"),
   879 => (x"7a",x"69",x"73",x"52"),
   880 => (x"25",x"20",x"3a",x"65"),
   881 => (x"70",x"20",x"2c",x"64"),
   882 => (x"69",x"74",x"72",x"61"),
   883 => (x"6e",x"6f",x"69",x"74"),
   884 => (x"65",x"7a",x"69",x"73"),
   885 => (x"64",x"25",x"20",x"3a"),
   886 => (x"66",x"6f",x"20",x"2c"),
   887 => (x"74",x"65",x"73",x"66"),
   888 => (x"20",x"66",x"6f",x"20"),
   889 => (x"3a",x"67",x"69",x"73"),
   890 => (x"2c",x"64",x"25",x"20"),
   891 => (x"67",x"69",x"73",x"20"),
   892 => (x"25",x"78",x"30",x"20"),
   893 => (x"52",x"00",x"0a",x"78"),
   894 => (x"69",x"64",x"61",x"65"),
   895 => (x"62",x"20",x"67",x"6e"),
   896 => (x"20",x"74",x"6f",x"6f"),
   897 => (x"74",x"63",x"65",x"73"),
   898 => (x"25",x"20",x"72",x"6f"),
   899 => (x"52",x"00",x"0a",x"64"),
   900 => (x"20",x"64",x"61",x"65"),
   901 => (x"74",x"6f",x"6f",x"62"),
   902 => (x"63",x"65",x"73",x"20"),
   903 => (x"20",x"72",x"6f",x"74"),
   904 => (x"6d",x"6f",x"72",x"66"),
   905 => (x"72",x"69",x"66",x"20"),
   906 => (x"70",x"20",x"74",x"73"),
   907 => (x"69",x"74",x"72",x"61"),
   908 => (x"6e",x"6f",x"69",x"74"),
   909 => (x"6e",x"55",x"00",x"0a"),
   910 => (x"70",x"70",x"75",x"73"),
   911 => (x"65",x"74",x"72",x"6f"),
   912 => (x"61",x"70",x"20",x"64"),
   913 => (x"74",x"69",x"74",x"72"),
   914 => (x"20",x"6e",x"6f",x"69"),
   915 => (x"65",x"70",x"79",x"74"),
   916 => (x"46",x"00",x"0d",x"21"),
   917 => (x"32",x"33",x"54",x"41"),
   918 => (x"00",x"20",x"20",x"20"),
   919 => (x"64",x"61",x"65",x"52"),
   920 => (x"20",x"67",x"6e",x"69"),
   921 => (x"0a",x"52",x"42",x"4d"),
   922 => (x"52",x"42",x"4d",x"00"),
   923 => (x"63",x"75",x"73",x"20"),
   924 => (x"73",x"73",x"65",x"63"),
   925 => (x"6c",x"6c",x"75",x"66"),
   926 => (x"65",x"72",x"20",x"79"),
   927 => (x"00",x"0a",x"64",x"61"),
   928 => (x"31",x"54",x"41",x"46"),
   929 => (x"20",x"20",x"20",x"36"),
   930 => (x"54",x"41",x"46",x"00"),
   931 => (x"20",x"20",x"32",x"33"),
   932 => (x"61",x"50",x"00",x"20"),
   933 => (x"74",x"69",x"74",x"72"),
   934 => (x"63",x"6e",x"6f",x"69"),
   935 => (x"74",x"6e",x"75",x"6f"),
   936 => (x"0a",x"64",x"25",x"20"),
   937 => (x"6e",x"75",x"48",x"00"),
   938 => (x"67",x"6e",x"69",x"74"),
   939 => (x"72",x"6f",x"66",x"20"),
   940 => (x"6c",x"69",x"66",x"20"),
   941 => (x"73",x"79",x"73",x"65"),
   942 => (x"0a",x"6d",x"65",x"74"),
   943 => (x"54",x"41",x"46",x"00"),
   944 => (x"20",x"20",x"32",x"33"),
   945 => (x"41",x"46",x"00",x"20"),
   946 => (x"20",x"36",x"31",x"54"),
   947 => (x"43",x"00",x"20",x"20"),
   948 => (x"74",x"73",x"75",x"6c"),
   949 => (x"73",x"20",x"72",x"65"),
   950 => (x"3a",x"65",x"7a",x"69"),
   951 => (x"2c",x"64",x"25",x"20"),
   952 => (x"75",x"6c",x"43",x"20"),
   953 => (x"72",x"65",x"74",x"73"),
   954 => (x"73",x"61",x"6d",x"20"),
   955 => (x"25",x"20",x"2c",x"6b"),
   956 => (x"0e",x"00",x"0a",x"64"),
   957 => (x"5d",x"5c",x"5b",x"5e"),
   958 => (x"c1",x"4a",x"71",x"0e"),
   959 => (x"02",x"bf",x"c2",x"eb"),
   960 => (x"4d",x"72",x"87",x"cc"),
   961 => (x"72",x"2d",x"b7",x"c7"),
   962 => (x"9b",x"ff",x"c1",x"4b"),
   963 => (x"4d",x"72",x"87",x"ca"),
   964 => (x"72",x"2d",x"b7",x"c8"),
   965 => (x"9b",x"ff",x"c3",x"4b"),
   966 => (x"1e",x"fa",x"e2",x"c1"),
   967 => (x"eb",x"c1",x"4a",x"75"),
   968 => (x"72",x"82",x"bf",x"c6"),
   969 => (x"87",x"f7",x"e3",x"49"),
   970 => (x"98",x"70",x"86",x"c4"),
   971 => (x"c0",x"87",x"c5",x"05"),
   972 => (x"87",x"e6",x"c0",x"48"),
   973 => (x"bf",x"c2",x"eb",x"c1"),
   974 => (x"73",x"87",x"d2",x"02"),
   975 => (x"c1",x"91",x"c4",x"49"),
   976 => (x"69",x"81",x"fa",x"e2"),
   977 => (x"ff",x"ff",x"cf",x"4c"),
   978 => (x"cb",x"9c",x"ff",x"ff"),
   979 => (x"c2",x"49",x"73",x"87"),
   980 => (x"fa",x"e2",x"c1",x"91"),
   981 => (x"4c",x"69",x"9f",x"81"),
   982 => (x"de",x"ec",x"48",x"74"),
   983 => (x"5b",x"5e",x"0e",x"87"),
   984 => (x"f4",x"0e",x"5d",x"5c"),
   985 => (x"c0",x"4c",x"71",x"86"),
   986 => (x"ce",x"eb",x"c1",x"4b"),
   987 => (x"eb",x"c1",x"4d",x"bf"),
   988 => (x"c1",x"7e",x"bf",x"d2"),
   989 => (x"02",x"bf",x"c2",x"eb"),
   990 => (x"ea",x"c1",x"87",x"c9"),
   991 => (x"c4",x"4a",x"bf",x"fa"),
   992 => (x"c1",x"87",x"c7",x"32"),
   993 => (x"4a",x"bf",x"d6",x"eb"),
   994 => (x"a6",x"c8",x"32",x"c4"),
   995 => (x"48",x"a6",x"c8",x"5a"),
   996 => (x"66",x"c4",x"78",x"c0"),
   997 => (x"06",x"a8",x"c0",x"48"),
   998 => (x"c8",x"87",x"e7",x"c2"),
   999 => (x"99",x"cf",x"49",x"66"),
  1000 => (x"c1",x"87",x"db",x"05"),
  1001 => (x"c4",x"1e",x"fa",x"e2"),
  1002 => (x"66",x"c4",x"49",x"66"),
  1003 => (x"c8",x"80",x"c1",x"48"),
  1004 => (x"e1",x"71",x"58",x"a6"),
  1005 => (x"86",x"c4",x"87",x"e9"),
  1006 => (x"4b",x"fa",x"e2",x"c1"),
  1007 => (x"e0",x"c0",x"87",x"c3"),
  1008 => (x"49",x"6b",x"97",x"83"),
  1009 => (x"ea",x"c1",x"02",x"99"),
  1010 => (x"49",x"6b",x"97",x"87"),
  1011 => (x"02",x"a9",x"e5",x"c3"),
  1012 => (x"cb",x"87",x"e0",x"c1"),
  1013 => (x"69",x"97",x"49",x"a3"),
  1014 => (x"05",x"99",x"d8",x"49"),
  1015 => (x"73",x"87",x"d4",x"c1"),
  1016 => (x"c3",x"ce",x"ff",x"49"),
  1017 => (x"c0",x"1e",x"cb",x"87"),
  1018 => (x"73",x"1e",x"66",x"e0"),
  1019 => (x"87",x"c9",x"e9",x"49"),
  1020 => (x"98",x"70",x"86",x"c8"),
  1021 => (x"87",x"fb",x"c0",x"05"),
  1022 => (x"c4",x"4a",x"a3",x"dc"),
  1023 => (x"79",x"6a",x"49",x"a4"),
  1024 => (x"c8",x"4a",x"a3",x"da"),
  1025 => (x"6a",x"9f",x"49",x"a4"),
  1026 => (x"c1",x"7e",x"71",x"79"),
  1027 => (x"02",x"bf",x"c2",x"eb"),
  1028 => (x"a3",x"d4",x"87",x"cf"),
  1029 => (x"49",x"69",x"9f",x"49"),
  1030 => (x"ff",x"ff",x"c0",x"4a"),
  1031 => (x"c2",x"32",x"d0",x"9a"),
  1032 => (x"72",x"4a",x"c0",x"87"),
  1033 => (x"bf",x"6e",x"48",x"49"),
  1034 => (x"78",x"08",x"6e",x"80"),
  1035 => (x"48",x"c1",x"7c",x"c0"),
  1036 => (x"c8",x"87",x"c1",x"c1"),
  1037 => (x"80",x"c1",x"48",x"66"),
  1038 => (x"c4",x"58",x"a6",x"cc"),
  1039 => (x"fd",x"04",x"a8",x"66"),
  1040 => (x"eb",x"c1",x"87",x"d9"),
  1041 => (x"c0",x"02",x"bf",x"c2"),
  1042 => (x"49",x"75",x"87",x"e8"),
  1043 => (x"70",x"87",x"e4",x"fa"),
  1044 => (x"cf",x"49",x"4d",x"49"),
  1045 => (x"f8",x"ff",x"ff",x"ff"),
  1046 => (x"d5",x"02",x"a9",x"99"),
  1047 => (x"c2",x"49",x"75",x"87"),
  1048 => (x"fa",x"ea",x"c1",x"89"),
  1049 => (x"eb",x"c1",x"91",x"bf"),
  1050 => (x"71",x"48",x"bf",x"ca"),
  1051 => (x"fc",x"7e",x"70",x"80"),
  1052 => (x"48",x"c0",x"87",x"db"),
  1053 => (x"c2",x"e8",x"8e",x"f4"),
  1054 => (x"1e",x"73",x"1e",x"87"),
  1055 => (x"49",x"6a",x"4a",x"71"),
  1056 => (x"7a",x"71",x"81",x"c1"),
  1057 => (x"bf",x"fe",x"ea",x"c1"),
  1058 => (x"87",x"cb",x"05",x"99"),
  1059 => (x"6b",x"4b",x"a2",x"c8"),
  1060 => (x"87",x"df",x"f9",x"49"),
  1061 => (x"c1",x"7b",x"49",x"70"),
  1062 => (x"87",x"e3",x"e7",x"48"),
  1063 => (x"71",x"1e",x"73",x"1e"),
  1064 => (x"ca",x"eb",x"c1",x"4b"),
  1065 => (x"a3",x"c8",x"4a",x"bf"),
  1066 => (x"c2",x"49",x"69",x"49"),
  1067 => (x"fa",x"ea",x"c1",x"89"),
  1068 => (x"a2",x"71",x"91",x"bf"),
  1069 => (x"fe",x"ea",x"c1",x"4a"),
  1070 => (x"99",x"6b",x"49",x"bf"),
  1071 => (x"c8",x"4a",x"a2",x"71"),
  1072 => (x"49",x"72",x"1e",x"66"),
  1073 => (x"87",x"d7",x"dd",x"ff"),
  1074 => (x"98",x"70",x"86",x"c4"),
  1075 => (x"c0",x"87",x"c4",x"05"),
  1076 => (x"c1",x"87",x"c2",x"48"),
  1077 => (x"87",x"e7",x"e6",x"48"),
  1078 => (x"71",x"1e",x"73",x"1e"),
  1079 => (x"29",x"d8",x"49",x"4b"),
  1080 => (x"73",x"99",x"ff",x"c3"),
  1081 => (x"cf",x"2a",x"c8",x"4a"),
  1082 => (x"72",x"9a",x"c0",x"fc"),
  1083 => (x"c8",x"4a",x"73",x"b1"),
  1084 => (x"f0",x"ff",x"c0",x"32"),
  1085 => (x"72",x"9a",x"c0",x"c0"),
  1086 => (x"d8",x"4a",x"73",x"b1"),
  1087 => (x"c0",x"c0",x"ff",x"32"),
  1088 => (x"72",x"9a",x"c0",x"c0"),
  1089 => (x"c4",x"48",x"71",x"b1"),
  1090 => (x"26",x"4d",x"26",x"87"),
  1091 => (x"26",x"4b",x"26",x"4c"),
  1092 => (x"4f",x"4f",x"00",x"4f"),
  1093 => (x"1e",x"1e",x"73",x"1e"),
  1094 => (x"49",x"4a",x"bf",x"e0"),
  1095 => (x"99",x"c0",x"e0",x"c0"),
  1096 => (x"87",x"d4",x"c2",x"02"),
  1097 => (x"c3",x"9a",x"ff",x"c3"),
  1098 => (x"c9",x"05",x"aa",x"f0"),
  1099 => (x"c8",x"c7",x"c1",x"87"),
  1100 => (x"c1",x"78",x"c1",x"48"),
  1101 => (x"e0",x"c3",x"87",x"f6"),
  1102 => (x"87",x"c9",x"05",x"aa"),
  1103 => (x"48",x"cc",x"c7",x"c1"),
  1104 => (x"e7",x"c1",x"78",x"c1"),
  1105 => (x"aa",x"fa",x"c3",x"87"),
  1106 => (x"87",x"e0",x"c1",x"02"),
  1107 => (x"bf",x"cc",x"c7",x"c1"),
  1108 => (x"c2",x"87",x"c6",x"02"),
  1109 => (x"c2",x"49",x"a2",x"c0"),
  1110 => (x"71",x"49",x"72",x"87"),
  1111 => (x"c8",x"c7",x"c1",x"4b"),
  1112 => (x"e0",x"c0",x"02",x"bf"),
  1113 => (x"c4",x"49",x"73",x"87"),
  1114 => (x"c1",x"91",x"29",x"b7"),
  1115 => (x"73",x"81",x"f1",x"ca"),
  1116 => (x"c2",x"9a",x"cf",x"4a"),
  1117 => (x"72",x"48",x"c1",x"92"),
  1118 => (x"ff",x"4a",x"70",x"30"),
  1119 => (x"69",x"48",x"72",x"ba"),
  1120 => (x"db",x"79",x"70",x"98"),
  1121 => (x"c4",x"49",x"73",x"87"),
  1122 => (x"c1",x"91",x"29",x"b7"),
  1123 => (x"73",x"81",x"f1",x"ca"),
  1124 => (x"c2",x"9a",x"cf",x"4a"),
  1125 => (x"72",x"48",x"c3",x"92"),
  1126 => (x"48",x"4a",x"70",x"30"),
  1127 => (x"79",x"70",x"b0",x"69"),
  1128 => (x"48",x"cc",x"c7",x"c1"),
  1129 => (x"c7",x"c1",x"78",x"c0"),
  1130 => (x"78",x"c0",x"48",x"c8"),
  1131 => (x"49",x"4a",x"bf",x"e0"),
  1132 => (x"99",x"c0",x"e0",x"c0"),
  1133 => (x"87",x"ec",x"fd",x"05"),
  1134 => (x"70",x"87",x"f6",x"c4"),
  1135 => (x"87",x"c4",x"26",x"7e"),
  1136 => (x"4c",x"26",x"4d",x"26"),
  1137 => (x"4f",x"26",x"4b",x"26"),
  1138 => (x"00",x"00",x"00",x"00"),
  1139 => (x"00",x"00",x"00",x"00"),
  1140 => (x"f2",x"c7",x"c1",x"1e"),
  1141 => (x"cf",x"c6",x"ff",x"49"),
  1142 => (x"72",x"4a",x"c0",x"87"),
  1143 => (x"c1",x"91",x"c4",x"49"),
  1144 => (x"c0",x"81",x"f1",x"ca"),
  1145 => (x"d0",x"82",x"c1",x"79"),
  1146 => (x"ee",x"04",x"aa",x"b7"),
  1147 => (x"87",x"cb",x"c4",x"87"),
  1148 => (x"65",x"4b",x"4f",x"26"),
  1149 => (x"61",x"6f",x"62",x"79"),
  1150 => (x"69",x"20",x"64",x"72"),
  1151 => (x"20",x"74",x"69",x"6e"),
  1152 => (x"63",x"6e",x"75",x"66"),
  1153 => (x"6e",x"6f",x"69",x"74"),
  1154 => (x"73",x"1e",x"00",x"0a"),
  1155 => (x"49",x"4b",x"71",x"1e"),
  1156 => (x"91",x"29",x"b7",x"c4"),
  1157 => (x"81",x"f1",x"ca",x"c1"),
  1158 => (x"9a",x"cf",x"4a",x"73"),
  1159 => (x"48",x"c2",x"92",x"c2"),
  1160 => (x"4a",x"70",x"30",x"72"),
  1161 => (x"48",x"72",x"ba",x"ff"),
  1162 => (x"79",x"70",x"98",x"69"),
  1163 => (x"0e",x"87",x"d5",x"fe"),
  1164 => (x"0e",x"5c",x"5b",x"5e"),
  1165 => (x"c4",x"4a",x"4c",x"71"),
  1166 => (x"c1",x"92",x"2a",x"b7"),
  1167 => (x"74",x"82",x"f1",x"ca"),
  1168 => (x"c2",x"9b",x"cf",x"4b"),
  1169 => (x"73",x"49",x"6a",x"93"),
  1170 => (x"c2",x"99",x"c3",x"29"),
  1171 => (x"70",x"30",x"73",x"48"),
  1172 => (x"73",x"bb",x"ff",x"4b"),
  1173 => (x"70",x"98",x"6a",x"48"),
  1174 => (x"fd",x"48",x"71",x"7a"),
  1175 => (x"5e",x"0e",x"87",x"e4"),
  1176 => (x"71",x"0e",x"5c",x"5b"),
  1177 => (x"b7",x"c4",x"4a",x"4b"),
  1178 => (x"ca",x"c1",x"92",x"2a"),
  1179 => (x"49",x"73",x"82",x"f1"),
  1180 => (x"91",x"c2",x"99",x"cf"),
  1181 => (x"28",x"71",x"48",x"6a"),
  1182 => (x"99",x"c3",x"49",x"70"),
  1183 => (x"ac",x"c2",x"4c",x"71"),
  1184 => (x"73",x"87",x"de",x"05"),
  1185 => (x"29",x"b7",x"c4",x"49"),
  1186 => (x"f1",x"ca",x"c1",x"91"),
  1187 => (x"cf",x"4a",x"73",x"81"),
  1188 => (x"c2",x"92",x"c2",x"9a"),
  1189 => (x"70",x"30",x"72",x"48"),
  1190 => (x"72",x"ba",x"ff",x"4a"),
  1191 => (x"70",x"98",x"69",x"48"),
  1192 => (x"02",x"ac",x"c2",x"79"),
  1193 => (x"49",x"c0",x"87",x"c4"),
  1194 => (x"49",x"c1",x"87",x"c2"),
  1195 => (x"d1",x"fc",x"48",x"71"),
  1196 => (x"00",x"00",x"00",x"87"),
  1197 => (x"00",x"00",x"00",x"00"),
  1198 => (x"00",x"00",x"00",x"00"),
  1199 => (x"00",x"00",x"00",x"00"),
  1200 => (x"00",x"00",x"00",x"00"),
  1201 => (x"00",x"00",x"00",x"00"),
  1202 => (x"00",x"00",x"00",x"00"),
  1203 => (x"00",x"00",x"00",x"00"),
  1204 => (x"00",x"00",x"00",x"00"),
  1205 => (x"00",x"00",x"00",x"00"),
  1206 => (x"00",x"00",x"00",x"00"),
  1207 => (x"00",x"00",x"00",x"00"),
  1208 => (x"00",x"00",x"00",x"00"),
  1209 => (x"00",x"00",x"00",x"00"),
  1210 => (x"00",x"00",x"00",x"00"),
  1211 => (x"00",x"00",x"00",x"00"),
  1212 => (x"fe",x"1e",x"1e",x"00"),
  1213 => (x"48",x"7e",x"bf",x"f0"),
  1214 => (x"1e",x"4f",x"26",x"26"),
  1215 => (x"c1",x"48",x"f0",x"fe"),
  1216 => (x"1e",x"4f",x"26",x"78"),
  1217 => (x"bf",x"fd",x"d0",x"c1"),
  1218 => (x"c1",x"31",x"cb",x"49"),
  1219 => (x"4a",x"bf",x"f9",x"d0"),
  1220 => (x"b1",x"72",x"32",x"c8"),
  1221 => (x"4f",x"26",x"48",x"71"),
  1222 => (x"48",x"c0",x"f8",x"1e"),
  1223 => (x"d0",x"c1",x"78",x"71"),
  1224 => (x"78",x"c0",x"48",x"f1"),
  1225 => (x"71",x"1e",x"4f",x"26"),
  1226 => (x"f5",x"d0",x"c1",x"4a"),
  1227 => (x"c1",x"78",x"c0",x"48"),
  1228 => (x"c0",x"5a",x"f5",x"d0"),
  1229 => (x"26",x"87",x"c2",x"49"),
  1230 => (x"5b",x"5e",x"0e",x"4f"),
  1231 => (x"1e",x"0e",x"5d",x"5c"),
  1232 => (x"4c",x"c0",x"4a",x"71"),
  1233 => (x"c1",x"7e",x"ff",x"c0"),
  1234 => (x"aa",x"bf",x"f5",x"d0"),
  1235 => (x"87",x"d3",x"c1",x"02"),
  1236 => (x"99",x"c1",x"49",x"72"),
  1237 => (x"c1",x"87",x"cb",x"02"),
  1238 => (x"48",x"bf",x"f1",x"d0"),
  1239 => (x"d0",x"c1",x"88",x"c1"),
  1240 => (x"49",x"72",x"58",x"f5"),
  1241 => (x"cb",x"02",x"99",x"c2"),
  1242 => (x"f1",x"d0",x"c1",x"87"),
  1243 => (x"80",x"c1",x"48",x"bf"),
  1244 => (x"58",x"f5",x"d0",x"c1"),
  1245 => (x"bf",x"f1",x"d0",x"c1"),
  1246 => (x"a8",x"b7",x"c0",x"48"),
  1247 => (x"c1",x"87",x"c6",x"03"),
  1248 => (x"c1",x"48",x"f1",x"d0"),
  1249 => (x"f1",x"d0",x"c1",x"78"),
  1250 => (x"b7",x"c1",x"48",x"bf"),
  1251 => (x"87",x"c6",x"06",x"a8"),
  1252 => (x"48",x"f1",x"d0",x"c1"),
  1253 => (x"49",x"72",x"78",x"c0"),
  1254 => (x"c2",x"02",x"99",x"d0"),
  1255 => (x"c1",x"4c",x"c1",x"87"),
  1256 => (x"c1",x"5a",x"f9",x"d0"),
  1257 => (x"49",x"bf",x"f1",x"d0"),
  1258 => (x"87",x"cd",x"02",x"99"),
  1259 => (x"db",x"02",x"89",x"c1"),
  1260 => (x"c0",x"02",x"89",x"87"),
  1261 => (x"e9",x"c0",x"87",x"ec"),
  1262 => (x"f9",x"d0",x"c1",x"87"),
  1263 => (x"81",x"74",x"49",x"bf"),
  1264 => (x"d0",x"c1",x"99",x"c3"),
  1265 => (x"4b",x"71",x"59",x"fd"),
  1266 => (x"87",x"dd",x"93",x"c5"),
  1267 => (x"d0",x"c1",x"4b",x"d4"),
  1268 => (x"74",x"49",x"bf",x"fd"),
  1269 => (x"c1",x"d1",x"c1",x"b9"),
  1270 => (x"05",x"99",x"71",x"59"),
  1271 => (x"7e",x"d7",x"87",x"cb"),
  1272 => (x"d0",x"c1",x"87",x"c7"),
  1273 => (x"c5",x"4b",x"bf",x"f1"),
  1274 => (x"48",x"c4",x"f8",x"93"),
  1275 => (x"93",x"c3",x"78",x"6e"),
  1276 => (x"d1",x"c1",x"4d",x"c0"),
  1277 => (x"82",x"73",x"4a",x"c3"),
  1278 => (x"d0",x"4a",x"6a",x"97"),
  1279 => (x"c2",x"d1",x"c1",x"32"),
  1280 => (x"97",x"81",x"73",x"49"),
  1281 => (x"31",x"c8",x"49",x"69"),
  1282 => (x"d1",x"c1",x"b2",x"71"),
  1283 => (x"81",x"73",x"49",x"c1"),
  1284 => (x"b2",x"49",x"69",x"97"),
  1285 => (x"91",x"c4",x"49",x"75"),
  1286 => (x"72",x"81",x"c8",x"f8"),
  1287 => (x"c1",x"83",x"c3",x"79"),
  1288 => (x"ad",x"b7",x"c5",x"85"),
  1289 => (x"87",x"ca",x"ff",x"04"),
  1290 => (x"26",x"4d",x"26",x"26"),
  1291 => (x"26",x"4b",x"26",x"4c"),
  1292 => (x"00",x"00",x"00",x"4f"),
  1293 => (x"00",x"00",x"00",x"00"),
  1294 => (x"00",x"00",x"00",x"00"),
  1295 => (x"00",x"00",x"00",x"00"),
  1296 => (x"00",x"3b",x"db",x"00"),
  1297 => (x"d5",x"00",x"48",x"55"),
  1298 => (x"48",x"51",x"00",x"49"),
  1299 => (x"00",x"3b",x"d1",x"00"),
  1300 => (x"21",x"08",x"b8",x"cf"),
  1301 => (x"19",x"27",x"05",x"05"),
  1302 => (x"02",x"21",x"e1",x"02"),
  1303 => (x"c9",x"02",x"1d",x"2f"),
  1304 => (x"a5",x"29",x"03",x"9c"),
  1305 => (x"04",x"a5",x"2f",x"04"),
  1306 => (x"29",x"04",x"9d",x"e9"),
  1307 => (x"bc",x"ef",x"03",x"a5"),
  1308 => (x"00",x"85",x"21",x"07"),
  1309 => (x"e1",x"03",x"9d",x"27"),
  1310 => (x"bd",x"21",x"00",x"84"),
  1311 => (x"fb",x"3d",x"26",x"07"),
  1312 => (x"e1",x"24",x"85",x"29"),
  1313 => (x"85",x"29",x"24",x"9d"),
  1314 => (x"24",x"bd",x"26",x"27"),
  1315 => (x"91",x"01",x"cc",x"61"),
  1316 => (x"52",x"91",x"02",x"52"),
  1317 => (x"02",x"5e",x"91",x"02"),
  1318 => (x"ef",x"a9",x"d2",x"67"),
  1319 => (x"a5",x"21",x"73",x"1c"),
  1320 => (x"94",x"a5",x"27",x"94"),
  1321 => (x"2f",x"74",x"9c",x"e1"),
  1322 => (x"5e",x"0e",x"93",x"25"),
  1323 => (x"0e",x"5d",x"5c",x"5b"),
  1324 => (x"c0",x"86",x"d8",x"ff"),
  1325 => (x"48",x"a6",x"c4",x"7e"),
  1326 => (x"78",x"bf",x"c4",x"fd"),
  1327 => (x"49",x"e3",x"e1",x"c1"),
  1328 => (x"87",x"e4",x"fa",x"fe"),
  1329 => (x"87",x"f2",x"c7",x"ff"),
  1330 => (x"d0",x"02",x"98",x"70"),
  1331 => (x"f2",x"d6",x"ff",x"87"),
  1332 => (x"02",x"98",x"70",x"87"),
  1333 => (x"a6",x"c8",x"87",x"c7"),
  1334 => (x"c5",x"78",x"c1",x"48"),
  1335 => (x"48",x"a6",x"c8",x"87"),
  1336 => (x"66",x"c8",x"78",x"c0"),
  1337 => (x"87",x"e0",x"c2",x"02"),
  1338 => (x"1e",x"f9",x"e1",x"c1"),
  1339 => (x"49",x"ea",x"eb",x"c1"),
  1340 => (x"c4",x"87",x"ea",x"e9"),
  1341 => (x"02",x"98",x"70",x"86"),
  1342 => (x"c8",x"87",x"cd",x"c2"),
  1343 => (x"eb",x"c1",x"48",x"a6"),
  1344 => (x"c1",x"78",x"bf",x"ee"),
  1345 => (x"87",x"d0",x"f8",x"49"),
  1346 => (x"d9",x"f8",x"49",x"c5"),
  1347 => (x"e6",x"e0",x"c1",x"87"),
  1348 => (x"d3",x"f9",x"fe",x"49"),
  1349 => (x"c1",x"48",x"f8",x"87"),
  1350 => (x"02",x"66",x"c8",x"78"),
  1351 => (x"c8",x"87",x"d6",x"c1"),
  1352 => (x"e2",x"c1",x"4c",x"66"),
  1353 => (x"eb",x"c1",x"1e",x"fa"),
  1354 => (x"ef",x"ed",x"49",x"ea"),
  1355 => (x"70",x"86",x"c4",x"87"),
  1356 => (x"87",x"c5",x"05",x"98"),
  1357 => (x"e2",x"cb",x"48",x"c0"),
  1358 => (x"b7",x"c0",x"c8",x"87"),
  1359 => (x"87",x"c4",x"04",x"ac"),
  1360 => (x"87",x"c4",x"8c",x"4a"),
  1361 => (x"4c",x"c0",x"4a",x"74"),
  1362 => (x"4b",x"fa",x"e2",x"c1"),
  1363 => (x"8a",x"c1",x"49",x"72"),
  1364 => (x"d3",x"02",x"99",x"71"),
  1365 => (x"fe",x"48",x"13",x"87"),
  1366 => (x"fc",x"b8",x"80",x"c0"),
  1367 => (x"49",x"72",x"78",x"08"),
  1368 => (x"99",x"71",x"8a",x"c1"),
  1369 => (x"87",x"ed",x"ff",x"05"),
  1370 => (x"49",x"ea",x"eb",x"c1"),
  1371 => (x"74",x"87",x"ca",x"ec"),
  1372 => (x"ed",x"fe",x"05",x"9c"),
  1373 => (x"c0",x"48",x"f8",x"87"),
  1374 => (x"ff",x"e0",x"c1",x"78"),
  1375 => (x"e7",x"f7",x"fe",x"49"),
  1376 => (x"f6",x"49",x"c0",x"87"),
  1377 => (x"87",x"d8",x"87",x"d2"),
  1378 => (x"cb",x"f6",x"49",x"c1"),
  1379 => (x"f6",x"49",x"c6",x"87"),
  1380 => (x"e1",x"c1",x"87",x"d4"),
  1381 => (x"f7",x"fe",x"49",x"c5"),
  1382 => (x"f4",x"ed",x"87",x"ce"),
  1383 => (x"87",x"fa",x"ff",x"87"),
  1384 => (x"a6",x"c8",x"4b",x"c0"),
  1385 => (x"4c",x"78",x"c0",x"48"),
  1386 => (x"c4",x"fd",x"80",x"c4"),
  1387 => (x"d8",x"c1",x"78",x"bf"),
  1388 => (x"87",x"fb",x"f1",x"49"),
  1389 => (x"c0",x"02",x"98",x"70"),
  1390 => (x"e0",x"c0",x"87",x"c3"),
  1391 => (x"f1",x"49",x"d2",x"b4"),
  1392 => (x"98",x"70",x"87",x"ed"),
  1393 => (x"87",x"c2",x"c0",x"02"),
  1394 => (x"49",x"d4",x"b4",x"d0"),
  1395 => (x"70",x"87",x"e0",x"f1"),
  1396 => (x"c3",x"c0",x"02",x"98"),
  1397 => (x"b4",x"e0",x"c0",x"87"),
  1398 => (x"d2",x"f1",x"49",x"d1"),
  1399 => (x"02",x"98",x"70",x"87"),
  1400 => (x"d0",x"87",x"c2",x"c0"),
  1401 => (x"f1",x"49",x"dd",x"b4"),
  1402 => (x"98",x"70",x"87",x"c5"),
  1403 => (x"87",x"c2",x"c0",x"02"),
  1404 => (x"49",x"db",x"b4",x"c1"),
  1405 => (x"70",x"87",x"f8",x"f0"),
  1406 => (x"c2",x"c0",x"02",x"98"),
  1407 => (x"dc",x"b4",x"c2",x"87"),
  1408 => (x"87",x"eb",x"f0",x"49"),
  1409 => (x"c0",x"02",x"98",x"70"),
  1410 => (x"b4",x"c4",x"87",x"c2"),
  1411 => (x"f0",x"49",x"e3",x"c0"),
  1412 => (x"98",x"70",x"87",x"dd"),
  1413 => (x"87",x"c2",x"c0",x"02"),
  1414 => (x"da",x"c1",x"b4",x"c8"),
  1415 => (x"87",x"cf",x"f0",x"49"),
  1416 => (x"c0",x"02",x"98",x"70"),
  1417 => (x"b3",x"d0",x"87",x"c2"),
  1418 => (x"f0",x"49",x"d9",x"c1"),
  1419 => (x"98",x"70",x"87",x"c1"),
  1420 => (x"87",x"c3",x"c0",x"02"),
  1421 => (x"c2",x"b3",x"e0",x"c0"),
  1422 => (x"f2",x"ef",x"49",x"d4"),
  1423 => (x"02",x"98",x"70",x"87"),
  1424 => (x"d0",x"87",x"c2",x"c0"),
  1425 => (x"49",x"d1",x"c2",x"b3"),
  1426 => (x"70",x"87",x"e4",x"ef"),
  1427 => (x"c3",x"c0",x"02",x"98"),
  1428 => (x"b3",x"e0",x"c0",x"87"),
  1429 => (x"ef",x"49",x"f5",x"c3"),
  1430 => (x"98",x"70",x"87",x"d5"),
  1431 => (x"87",x"c2",x"c0",x"02"),
  1432 => (x"f2",x"c3",x"b3",x"c1"),
  1433 => (x"87",x"c7",x"ef",x"49"),
  1434 => (x"c0",x"02",x"98",x"70"),
  1435 => (x"b3",x"c2",x"87",x"c2"),
  1436 => (x"ee",x"49",x"eb",x"c3"),
  1437 => (x"98",x"70",x"87",x"f9"),
  1438 => (x"87",x"c2",x"c0",x"02"),
  1439 => (x"f4",x"c3",x"b3",x"c4"),
  1440 => (x"87",x"eb",x"ee",x"49"),
  1441 => (x"c0",x"02",x"98",x"70"),
  1442 => (x"b3",x"c8",x"87",x"c2"),
  1443 => (x"ee",x"49",x"f1",x"c0"),
  1444 => (x"98",x"70",x"87",x"dd"),
  1445 => (x"87",x"c8",x"c0",x"02"),
  1446 => (x"d0",x"48",x"66",x"c8"),
  1447 => (x"58",x"a6",x"cc",x"b0"),
  1448 => (x"ee",x"49",x"f2",x"c0"),
  1449 => (x"98",x"70",x"87",x"c9"),
  1450 => (x"87",x"c9",x"c0",x"02"),
  1451 => (x"c0",x"48",x"66",x"c8"),
  1452 => (x"a6",x"cc",x"b0",x"e0"),
  1453 => (x"49",x"c3",x"c1",x"58"),
  1454 => (x"70",x"87",x"f4",x"ed"),
  1455 => (x"c8",x"c0",x"02",x"98"),
  1456 => (x"48",x"66",x"c8",x"87"),
  1457 => (x"a6",x"cc",x"b0",x"c1"),
  1458 => (x"49",x"c2",x"c1",x"58"),
  1459 => (x"70",x"87",x"e0",x"ed"),
  1460 => (x"c8",x"c0",x"02",x"98"),
  1461 => (x"48",x"66",x"c8",x"87"),
  1462 => (x"a6",x"cc",x"b0",x"c2"),
  1463 => (x"49",x"fb",x"c0",x"58"),
  1464 => (x"70",x"87",x"cc",x"ed"),
  1465 => (x"c8",x"c0",x"02",x"98"),
  1466 => (x"48",x"66",x"c8",x"87"),
  1467 => (x"a6",x"cc",x"b0",x"c4"),
  1468 => (x"49",x"cb",x"c1",x"58"),
  1469 => (x"70",x"87",x"f8",x"ec"),
  1470 => (x"c8",x"c0",x"02",x"98"),
  1471 => (x"48",x"66",x"c8",x"87"),
  1472 => (x"a6",x"cc",x"b0",x"c8"),
  1473 => (x"4d",x"66",x"cc",x"58"),
  1474 => (x"ee",x"c0",x"9d",x"c1"),
  1475 => (x"87",x"df",x"ec",x"49"),
  1476 => (x"c0",x"02",x"98",x"70"),
  1477 => (x"b5",x"c1",x"87",x"c2"),
  1478 => (x"ec",x"49",x"f6",x"c0"),
  1479 => (x"98",x"70",x"87",x"d1"),
  1480 => (x"87",x"c2",x"c0",x"02"),
  1481 => (x"fd",x"c0",x"b5",x"c2"),
  1482 => (x"87",x"c3",x"ec",x"49"),
  1483 => (x"c0",x"02",x"98",x"70"),
  1484 => (x"b5",x"c4",x"87",x"c2"),
  1485 => (x"f6",x"eb",x"49",x"d6"),
  1486 => (x"02",x"98",x"70",x"87"),
  1487 => (x"c8",x"87",x"c2",x"c0"),
  1488 => (x"eb",x"49",x"de",x"b5"),
  1489 => (x"98",x"70",x"87",x"e9"),
  1490 => (x"87",x"c2",x"c0",x"02"),
  1491 => (x"e6",x"c0",x"b5",x"d0"),
  1492 => (x"87",x"db",x"eb",x"49"),
  1493 => (x"c0",x"02",x"98",x"70"),
  1494 => (x"e0",x"c0",x"87",x"c3"),
  1495 => (x"eb",x"49",x"c6",x"b5"),
  1496 => (x"98",x"70",x"87",x"cd"),
  1497 => (x"87",x"c3",x"c0",x"02"),
  1498 => (x"c7",x"b5",x"c0",x"c4"),
  1499 => (x"87",x"ee",x"eb",x"49"),
  1500 => (x"c0",x"05",x"98",x"70"),
  1501 => (x"66",x"cc",x"87",x"d2"),
  1502 => (x"02",x"99",x"d0",x"49"),
  1503 => (x"c4",x"87",x"f8",x"c0"),
  1504 => (x"99",x"d0",x"49",x"66"),
  1505 => (x"87",x"ef",x"c0",x"05"),
  1506 => (x"fd",x"e9",x"49",x"c7"),
  1507 => (x"c1",x"48",x"6e",x"87"),
  1508 => (x"49",x"7e",x"70",x"b8"),
  1509 => (x"6e",x"87",x"c1",x"ee"),
  1510 => (x"d5",x"e1",x"c1",x"1e"),
  1511 => (x"d9",x"ee",x"fe",x"1e"),
  1512 => (x"6e",x"86",x"c8",x"87"),
  1513 => (x"87",x"cf",x"c0",x"05"),
  1514 => (x"70",x"87",x"d8",x"ed"),
  1515 => (x"b2",x"c1",x"4a",x"49"),
  1516 => (x"78",x"72",x"48",x"f4"),
  1517 => (x"fd",x"78",x"71",x"78"),
  1518 => (x"78",x"75",x"48",x"c4"),
  1519 => (x"31",x"d0",x"49",x"73"),
  1520 => (x"c8",x"4a",x"66",x"c8"),
  1521 => (x"74",x"b1",x"72",x"32"),
  1522 => (x"48",x"c8",x"fd",x"b1"),
  1523 => (x"48",x"68",x"78",x"71"),
  1524 => (x"c8",x"98",x"ff",x"c0"),
  1525 => (x"a6",x"d4",x"58",x"a6"),
  1526 => (x"48",x"66",x"d0",x"5b"),
  1527 => (x"d8",x"b0",x"66",x"c4"),
  1528 => (x"4b",x"70",x"58",x"a6"),
  1529 => (x"48",x"bf",x"c8",x"fd"),
  1530 => (x"a6",x"dc",x"28",x"c8"),
  1531 => (x"98",x"ff",x"c0",x"58"),
  1532 => (x"58",x"a6",x"e0",x"c0"),
  1533 => (x"5b",x"a6",x"e4",x"c0"),
  1534 => (x"48",x"66",x"e0",x"c0"),
  1535 => (x"c0",x"b0",x"66",x"dc"),
  1536 => (x"70",x"58",x"a6",x"e8"),
  1537 => (x"c0",x"02",x"6e",x"4b"),
  1538 => (x"49",x"73",x"87",x"c5"),
  1539 => (x"c4",x"87",x"ea",x"ec"),
  1540 => (x"66",x"cc",x"48",x"a6"),
  1541 => (x"87",x"fc",x"e3",x"78"),
  1542 => (x"ff",x"87",x"c5",x"f6"),
  1543 => (x"4d",x"26",x"8e",x"d8"),
  1544 => (x"4b",x"26",x"4c",x"26"),
  1545 => (x"70",x"4f",x"4f",x"26"),
  1546 => (x"64",x"65",x"6e",x"65"),
  1547 => (x"6c",x"69",x"66",x"20"),
  1548 => (x"6c",x"20",x"2c",x"65"),
  1549 => (x"69",x"64",x"61",x"6f"),
  1550 => (x"2e",x"2e",x"67",x"6e"),
  1551 => (x"44",x"00",x"0a",x"2e"),
  1552 => (x"0a",x"65",x"6e",x"6f"),
  1553 => (x"20",x"44",x"53",x"00"),
  1554 => (x"74",x"6f",x"6f",x"62"),
  1555 => (x"69",x"61",x"66",x"20"),
  1556 => (x"0a",x"64",x"65",x"6c"),
  1557 => (x"6f",x"68",x"53",x"00"),
  1558 => (x"65",x"6d",x"20",x"77"),
  1559 => (x"25",x"20",x"75",x"6e"),
  1560 => (x"49",x"00",x"0a",x"64"),
  1561 => (x"69",x"74",x"69",x"6e"),
  1562 => (x"7a",x"69",x"6c",x"61"),
  1563 => (x"20",x"67",x"6e",x"69"),
  1564 => (x"63",x"20",x"44",x"53"),
  1565 => (x"0a",x"64",x"72",x"61"),
  1566 => (x"4d",x"41",x"52",x"00"),
  1567 => (x"45",x"47",x"41",x"50"),
  1568 => (x"4d",x"4f",x"52",x"20"),
  1569 => (x"00",x"11",x"d0",x"00"),
  1570 => (x"00",x"11",x"d0",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

