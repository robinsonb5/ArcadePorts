
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity Boot_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of Boot_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"2c",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"29"),
    10 => (x"87",x"fd",x"00",x"4f"),
    11 => (x"e4",x"ee",x"c1",x"4f"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"00",x"1b",x"a4",x"27"),
    14 => (x"20",x"27",x"49",x"00"),
    15 => (x"48",x"00",x"00",x"19"),
    16 => (x"c0",x"05",x"a9",x"70"),
    17 => (x"27",x"87",x"f9",x"50"),
    18 => (x"00",x"00",x"19",x"1d"),
    19 => (x"19",x"19",x"27",x"4c"),
    20 => (x"74",x"4d",x"00",x"00"),
    21 => (x"87",x"c6",x"02",x"ad"),
    22 => (x"0f",x"6c",x"8c",x"c4"),
    23 => (x"d3",x"c1",x"87",x"f5"),
    24 => (x"1d",x"27",x"87",x"eb"),
    25 => (x"4c",x"00",x"00",x"19"),
    26 => (x"00",x"19",x"1d",x"27"),
    27 => (x"ad",x"74",x"4d",x"00"),
    28 => (x"24",x"87",x"c4",x"02"),
    29 => (x"00",x"87",x"f7",x"0f"),
    30 => (x"1e",x"1e",x"87",x"fd"),
    31 => (x"69",x"49",x"c0",x"ff"),
    32 => (x"98",x"c0",x"c4",x"48"),
    33 => (x"6e",x"58",x"a6",x"c4"),
    34 => (x"c8",x"87",x"f4",x"02"),
    35 => (x"26",x"48",x"79",x"66"),
    36 => (x"4d",x"26",x"87",x"c6"),
    37 => (x"4b",x"26",x"4c",x"26"),
    38 => (x"5e",x"0e",x"4f",x"26"),
    39 => (x"cc",x"0e",x"5c",x"5b"),
    40 => (x"4b",x"c0",x"4c",x"66"),
    41 => (x"ff",x"c3",x"4a",x"14"),
    42 => (x"02",x"9a",x"72",x"9a"),
    43 => (x"49",x"72",x"87",x"d5"),
    44 => (x"c5",x"ff",x"1e",x"71"),
    45 => (x"c1",x"86",x"c4",x"87"),
    46 => (x"c3",x"4a",x"14",x"83"),
    47 => (x"9a",x"72",x"9a",x"ff"),
    48 => (x"73",x"87",x"eb",x"05"),
    49 => (x"87",x"cc",x"ff",x"48"),
    50 => (x"5c",x"5b",x"5e",x"0e"),
    51 => (x"86",x"f0",x"0e",x"5d"),
    52 => (x"a6",x"c4",x"4b",x"c0"),
    53 => (x"c0",x"78",x"c0",x"48"),
    54 => (x"c0",x"4c",x"a6",x"e4"),
    55 => (x"48",x"49",x"66",x"e0"),
    56 => (x"e4",x"c0",x"80",x"c1"),
    57 => (x"4a",x"11",x"58",x"a6"),
    58 => (x"ba",x"82",x"c0",x"fe"),
    59 => (x"c4",x"02",x"9a",x"72"),
    60 => (x"66",x"c4",x"87",x"d3"),
    61 => (x"87",x"e2",x"c3",x"02"),
    62 => (x"c0",x"48",x"a6",x"c4"),
    63 => (x"c0",x"49",x"72",x"78"),
    64 => (x"c2",x"02",x"aa",x"f0"),
    65 => (x"e3",x"c1",x"87",x"f2"),
    66 => (x"f3",x"c2",x"02",x"a9"),
    67 => (x"a9",x"e4",x"c1",x"87"),
    68 => (x"87",x"e1",x"c0",x"02"),
    69 => (x"02",x"a9",x"ec",x"c1"),
    70 => (x"c1",x"87",x"dd",x"c2"),
    71 => (x"d4",x"02",x"a9",x"f0"),
    72 => (x"a9",x"f3",x"c1",x"87"),
    73 => (x"87",x"fc",x"c1",x"02"),
    74 => (x"02",x"a9",x"f5",x"c1"),
    75 => (x"f8",x"c1",x"87",x"c7"),
    76 => (x"dc",x"c2",x"05",x"a9"),
    77 => (x"74",x"84",x"c4",x"87"),
    78 => (x"76",x"89",x"c4",x"49"),
    79 => (x"6e",x"78",x"69",x"48"),
    80 => (x"87",x"d3",x"c1",x"02"),
    81 => (x"78",x"c0",x"80",x"c8"),
    82 => (x"c0",x"48",x"a6",x"cc"),
    83 => (x"dc",x"49",x"6e",x"78"),
    84 => (x"4a",x"71",x"29",x"b7"),
    85 => (x"48",x"6e",x"9a",x"cf"),
    86 => (x"a6",x"c4",x"30",x"c4"),
    87 => (x"02",x"9a",x"72",x"58"),
    88 => (x"a6",x"c8",x"87",x"c5"),
    89 => (x"c9",x"78",x"c1",x"48"),
    90 => (x"87",x"c5",x"06",x"aa"),
    91 => (x"c3",x"82",x"f7",x"c0"),
    92 => (x"82",x"f0",x"c0",x"87"),
    93 => (x"c9",x"02",x"66",x"c8"),
    94 => (x"fb",x"1e",x"72",x"87"),
    95 => (x"86",x"c4",x"87",x"fc"),
    96 => (x"66",x"cc",x"83",x"c1"),
    97 => (x"d0",x"80",x"c1",x"48"),
    98 => (x"66",x"cc",x"58",x"a6"),
    99 => (x"a8",x"b7",x"c8",x"48"),
   100 => (x"87",x"f9",x"fe",x"04"),
   101 => (x"c0",x"87",x"d7",x"c1"),
   102 => (x"dd",x"fb",x"1e",x"f0"),
   103 => (x"c1",x"86",x"c4",x"87"),
   104 => (x"87",x"ca",x"c1",x"83"),
   105 => (x"49",x"74",x"84",x"c4"),
   106 => (x"1e",x"69",x"89",x"c4"),
   107 => (x"c4",x"87",x"eb",x"fb"),
   108 => (x"71",x"49",x"70",x"86"),
   109 => (x"87",x"f6",x"c0",x"83"),
   110 => (x"c1",x"48",x"a6",x"c4"),
   111 => (x"87",x"ee",x"c0",x"78"),
   112 => (x"49",x"74",x"84",x"c4"),
   113 => (x"1e",x"69",x"89",x"c4"),
   114 => (x"c4",x"87",x"ef",x"fa"),
   115 => (x"dd",x"83",x"c1",x"86"),
   116 => (x"fa",x"1e",x"72",x"87"),
   117 => (x"86",x"c4",x"87",x"e4"),
   118 => (x"e5",x"c0",x"87",x"d4"),
   119 => (x"87",x"c7",x"05",x"aa"),
   120 => (x"c1",x"48",x"a6",x"c4"),
   121 => (x"72",x"87",x"c7",x"78"),
   122 => (x"87",x"ce",x"fa",x"1e"),
   123 => (x"e0",x"c0",x"86",x"c4"),
   124 => (x"c1",x"48",x"49",x"66"),
   125 => (x"a6",x"e4",x"c0",x"80"),
   126 => (x"fe",x"4a",x"11",x"58"),
   127 => (x"72",x"ba",x"82",x"c0"),
   128 => (x"ed",x"fb",x"05",x"9a"),
   129 => (x"f0",x"48",x"73",x"87"),
   130 => (x"26",x"4d",x"26",x"8e"),
   131 => (x"26",x"4b",x"26",x"4c"),
   132 => (x"0e",x"5e",x"0e",x"4f"),
   133 => (x"d4",x"ff",x"86",x"e8"),
   134 => (x"7a",x"ff",x"c3",x"4a"),
   135 => (x"ff",x"c3",x"49",x"6a"),
   136 => (x"c8",x"48",x"6a",x"7a"),
   137 => (x"58",x"a6",x"c4",x"30"),
   138 => (x"6e",x"59",x"a6",x"c8"),
   139 => (x"7a",x"ff",x"c3",x"b1"),
   140 => (x"30",x"d0",x"48",x"6a"),
   141 => (x"d0",x"58",x"a6",x"cc"),
   142 => (x"66",x"c8",x"59",x"a6"),
   143 => (x"7a",x"ff",x"c3",x"b1"),
   144 => (x"30",x"d8",x"48",x"6a"),
   145 => (x"d8",x"58",x"a6",x"d4"),
   146 => (x"66",x"d0",x"59",x"a6"),
   147 => (x"e8",x"48",x"71",x"b1"),
   148 => (x"26",x"87",x"c6",x"8e"),
   149 => (x"26",x"4c",x"26",x"4d"),
   150 => (x"0e",x"4f",x"26",x"4b"),
   151 => (x"86",x"f4",x"0e",x"5e"),
   152 => (x"c3",x"4a",x"d4",x"ff"),
   153 => (x"49",x"6a",x"7a",x"ff"),
   154 => (x"71",x"7a",x"ff",x"c3"),
   155 => (x"c4",x"30",x"c8",x"48"),
   156 => (x"49",x"6a",x"58",x"a6"),
   157 => (x"ff",x"c3",x"b1",x"6e"),
   158 => (x"c8",x"48",x"71",x"7a"),
   159 => (x"58",x"a6",x"c8",x"30"),
   160 => (x"66",x"c4",x"49",x"6a"),
   161 => (x"7a",x"ff",x"c3",x"b1"),
   162 => (x"30",x"c8",x"48",x"71"),
   163 => (x"6a",x"58",x"a6",x"cc"),
   164 => (x"b1",x"66",x"c8",x"49"),
   165 => (x"8e",x"f4",x"48",x"71"),
   166 => (x"0e",x"87",x"fe",x"fe"),
   167 => (x"0e",x"5c",x"5b",x"5e"),
   168 => (x"cc",x"4c",x"d4",x"ff"),
   169 => (x"ff",x"c3",x"48",x"66"),
   170 => (x"c1",x"7c",x"70",x"98"),
   171 => (x"05",x"bf",x"e4",x"e4"),
   172 => (x"66",x"d0",x"87",x"c8"),
   173 => (x"d4",x"30",x"c9",x"48"),
   174 => (x"66",x"d0",x"58",x"a6"),
   175 => (x"71",x"29",x"d8",x"49"),
   176 => (x"98",x"ff",x"c3",x"48"),
   177 => (x"66",x"d0",x"7c",x"70"),
   178 => (x"71",x"29",x"d0",x"49"),
   179 => (x"98",x"ff",x"c3",x"48"),
   180 => (x"66",x"d0",x"7c",x"70"),
   181 => (x"71",x"29",x"c8",x"49"),
   182 => (x"98",x"ff",x"c3",x"48"),
   183 => (x"66",x"d0",x"7c",x"70"),
   184 => (x"98",x"ff",x"c3",x"48"),
   185 => (x"66",x"cc",x"7c",x"70"),
   186 => (x"71",x"29",x"d0",x"49"),
   187 => (x"98",x"ff",x"c3",x"48"),
   188 => (x"4a",x"6c",x"7c",x"70"),
   189 => (x"4b",x"ff",x"f0",x"c9"),
   190 => (x"05",x"aa",x"ff",x"c3"),
   191 => (x"ff",x"c3",x"87",x"d0"),
   192 => (x"c1",x"4a",x"6c",x"7c"),
   193 => (x"87",x"c6",x"02",x"8b"),
   194 => (x"02",x"aa",x"ff",x"c3"),
   195 => (x"48",x"72",x"87",x"f0"),
   196 => (x"1e",x"87",x"c2",x"fd"),
   197 => (x"d4",x"ff",x"49",x"c0"),
   198 => (x"78",x"ff",x"c3",x"48"),
   199 => (x"c8",x"c3",x"81",x"c1"),
   200 => (x"f1",x"04",x"a9",x"b7"),
   201 => (x"87",x"f1",x"fc",x"87"),
   202 => (x"0e",x"5b",x"5e",x"0e"),
   203 => (x"f8",x"c4",x"87",x"e5"),
   204 => (x"1e",x"c0",x"4b",x"df"),
   205 => (x"c1",x"f0",x"ff",x"c0"),
   206 => (x"de",x"fd",x"1e",x"f7"),
   207 => (x"c1",x"86",x"c8",x"87"),
   208 => (x"ea",x"c0",x"05",x"a8"),
   209 => (x"48",x"d4",x"ff",x"87"),
   210 => (x"c1",x"78",x"ff",x"c3"),
   211 => (x"c0",x"c0",x"c0",x"c0"),
   212 => (x"e1",x"c0",x"1e",x"c0"),
   213 => (x"1e",x"e9",x"c1",x"f0"),
   214 => (x"c8",x"87",x"c0",x"fd"),
   215 => (x"05",x"98",x"70",x"86"),
   216 => (x"d4",x"ff",x"87",x"ca"),
   217 => (x"78",x"ff",x"c3",x"48"),
   218 => (x"87",x"cb",x"48",x"c1"),
   219 => (x"c1",x"87",x"e4",x"fe"),
   220 => (x"fd",x"fe",x"05",x"8b"),
   221 => (x"fb",x"48",x"c0",x"87"),
   222 => (x"5e",x"0e",x"87",x"dd"),
   223 => (x"d4",x"ff",x"0e",x"5b"),
   224 => (x"78",x"ff",x"c3",x"48"),
   225 => (x"1e",x"fb",x"e5",x"c0"),
   226 => (x"c4",x"87",x"cf",x"f4"),
   227 => (x"c0",x"4b",x"d3",x"86"),
   228 => (x"f0",x"ff",x"c0",x"1e"),
   229 => (x"fc",x"1e",x"c1",x"c1"),
   230 => (x"86",x"c8",x"87",x"c1"),
   231 => (x"ca",x"05",x"98",x"70"),
   232 => (x"48",x"d4",x"ff",x"87"),
   233 => (x"c1",x"78",x"ff",x"c3"),
   234 => (x"fd",x"87",x"cb",x"48"),
   235 => (x"8b",x"c1",x"87",x"e5"),
   236 => (x"87",x"db",x"ff",x"05"),
   237 => (x"de",x"fa",x"48",x"c0"),
   238 => (x"5b",x"5e",x"0e",x"87"),
   239 => (x"ff",x"0e",x"5d",x"5c"),
   240 => (x"ce",x"fd",x"4d",x"d4"),
   241 => (x"1e",x"ea",x"c6",x"87"),
   242 => (x"c1",x"f0",x"e1",x"c0"),
   243 => (x"ca",x"fb",x"1e",x"c8"),
   244 => (x"70",x"86",x"c8",x"87"),
   245 => (x"d3",x"1e",x"73",x"4b"),
   246 => (x"eb",x"f3",x"1e",x"c0"),
   247 => (x"c1",x"86",x"c8",x"87"),
   248 => (x"87",x"c8",x"02",x"ab"),
   249 => (x"c0",x"87",x"d3",x"fe"),
   250 => (x"87",x"cf",x"c2",x"48"),
   251 => (x"70",x"87",x"ec",x"f9"),
   252 => (x"ff",x"ff",x"cf",x"49"),
   253 => (x"a9",x"ea",x"c6",x"99"),
   254 => (x"fd",x"87",x"c8",x"02"),
   255 => (x"48",x"c0",x"87",x"fc"),
   256 => (x"c3",x"87",x"f8",x"c1"),
   257 => (x"f1",x"c0",x"7d",x"ff"),
   258 => (x"87",x"dc",x"fc",x"4c"),
   259 => (x"c1",x"02",x"98",x"70"),
   260 => (x"1e",x"c0",x"87",x"d0"),
   261 => (x"c1",x"f0",x"ff",x"c0"),
   262 => (x"fe",x"f9",x"1e",x"fa"),
   263 => (x"70",x"86",x"c8",x"87"),
   264 => (x"05",x"9b",x"73",x"4b"),
   265 => (x"73",x"87",x"f1",x"c0"),
   266 => (x"1e",x"fe",x"d1",x"1e"),
   267 => (x"c8",x"87",x"d9",x"f2"),
   268 => (x"7d",x"ff",x"c3",x"86"),
   269 => (x"1e",x"73",x"4b",x"6d"),
   270 => (x"f2",x"1e",x"ca",x"d2"),
   271 => (x"86",x"c8",x"87",x"ca"),
   272 => (x"7d",x"7d",x"ff",x"c3"),
   273 => (x"49",x"73",x"7d",x"7d"),
   274 => (x"02",x"99",x"c0",x"c1"),
   275 => (x"48",x"c1",x"87",x"c5"),
   276 => (x"c0",x"87",x"e8",x"c0"),
   277 => (x"87",x"e3",x"c0",x"48"),
   278 => (x"d8",x"d2",x"1e",x"73"),
   279 => (x"87",x"e8",x"f1",x"1e"),
   280 => (x"ac",x"c2",x"86",x"c8"),
   281 => (x"d2",x"87",x"cc",x"05"),
   282 => (x"db",x"f1",x"1e",x"e4"),
   283 => (x"c0",x"86",x"c4",x"87"),
   284 => (x"c1",x"87",x"c8",x"48"),
   285 => (x"d0",x"fe",x"05",x"8c"),
   286 => (x"f7",x"48",x"c0",x"87"),
   287 => (x"4d",x"43",x"87",x"d5"),
   288 => (x"20",x"38",x"35",x"44"),
   289 => (x"20",x"0a",x"64",x"25"),
   290 => (x"4d",x"43",x"00",x"20"),
   291 => (x"5f",x"38",x"35",x"44"),
   292 => (x"64",x"25",x"20",x"32"),
   293 => (x"00",x"20",x"20",x"0a"),
   294 => (x"35",x"44",x"4d",x"43"),
   295 => (x"64",x"25",x"20",x"38"),
   296 => (x"00",x"20",x"20",x"0a"),
   297 => (x"43",x"48",x"44",x"53"),
   298 => (x"69",x"6e",x"49",x"20"),
   299 => (x"6c",x"61",x"69",x"74"),
   300 => (x"74",x"61",x"7a",x"69"),
   301 => (x"20",x"6e",x"6f",x"69"),
   302 => (x"6f",x"72",x"72",x"65"),
   303 => (x"00",x"0a",x"21",x"72"),
   304 => (x"5f",x"64",x"6d",x"63"),
   305 => (x"38",x"44",x"4d",x"43"),
   306 => (x"73",x"65",x"72",x"20"),
   307 => (x"73",x"6e",x"6f",x"70"),
   308 => (x"25",x"20",x"3a",x"65"),
   309 => (x"0e",x"00",x"0a",x"64"),
   310 => (x"5d",x"5c",x"5b",x"5e"),
   311 => (x"d0",x"ff",x"1e",x"0e"),
   312 => (x"c0",x"c0",x"c8",x"4d"),
   313 => (x"e4",x"e4",x"c1",x"4b"),
   314 => (x"d6",x"78",x"c1",x"48"),
   315 => (x"e9",x"ee",x"1e",x"fb"),
   316 => (x"c7",x"86",x"c4",x"87"),
   317 => (x"73",x"48",x"6d",x"4c"),
   318 => (x"58",x"a6",x"c4",x"98"),
   319 => (x"cc",x"c0",x"02",x"6e"),
   320 => (x"73",x"48",x"6d",x"87"),
   321 => (x"58",x"a6",x"c4",x"98"),
   322 => (x"f4",x"ff",x"05",x"6e"),
   323 => (x"f8",x"7d",x"c2",x"87"),
   324 => (x"48",x"6d",x"87",x"c1"),
   325 => (x"a6",x"c4",x"98",x"73"),
   326 => (x"c0",x"02",x"6e",x"58"),
   327 => (x"48",x"6d",x"87",x"cc"),
   328 => (x"a6",x"c4",x"98",x"73"),
   329 => (x"ff",x"05",x"6e",x"58"),
   330 => (x"7d",x"c3",x"87",x"f4"),
   331 => (x"e5",x"c0",x"1e",x"c0"),
   332 => (x"1e",x"c0",x"c1",x"d0"),
   333 => (x"c8",x"87",x"e4",x"f5"),
   334 => (x"05",x"a8",x"c1",x"86"),
   335 => (x"c1",x"87",x"c2",x"c0"),
   336 => (x"05",x"ac",x"c2",x"4c"),
   337 => (x"d6",x"87",x"cd",x"c0"),
   338 => (x"cd",x"ed",x"1e",x"f6"),
   339 => (x"c0",x"86",x"c4",x"87"),
   340 => (x"87",x"de",x"c1",x"48"),
   341 => (x"fe",x"05",x"8c",x"c1"),
   342 => (x"dc",x"f9",x"87",x"db"),
   343 => (x"e8",x"e4",x"c1",x"87"),
   344 => (x"e4",x"e4",x"c1",x"58"),
   345 => (x"cd",x"c0",x"05",x"bf"),
   346 => (x"c0",x"1e",x"c1",x"87"),
   347 => (x"d0",x"c1",x"f0",x"ff"),
   348 => (x"87",x"e7",x"f4",x"1e"),
   349 => (x"d4",x"ff",x"86",x"c8"),
   350 => (x"78",x"ff",x"c3",x"48"),
   351 => (x"c1",x"87",x"c1",x"ca"),
   352 => (x"c1",x"58",x"ec",x"e4"),
   353 => (x"1e",x"bf",x"e8",x"e4"),
   354 => (x"ec",x"1e",x"ff",x"d6"),
   355 => (x"86",x"c8",x"87",x"fa"),
   356 => (x"98",x"73",x"48",x"6d"),
   357 => (x"6e",x"58",x"a6",x"c4"),
   358 => (x"87",x"cc",x"c0",x"02"),
   359 => (x"98",x"73",x"48",x"6d"),
   360 => (x"6e",x"58",x"a6",x"c4"),
   361 => (x"87",x"f4",x"ff",x"05"),
   362 => (x"d4",x"ff",x"7d",x"c2"),
   363 => (x"78",x"ff",x"c3",x"48"),
   364 => (x"f2",x"26",x"48",x"c1"),
   365 => (x"45",x"49",x"87",x"dd"),
   366 => (x"53",x"00",x"52",x"52"),
   367 => (x"53",x"00",x"49",x"50"),
   368 => (x"61",x"63",x"20",x"44"),
   369 => (x"73",x"20",x"64",x"72"),
   370 => (x"20",x"65",x"7a",x"69"),
   371 => (x"25",x"20",x"73",x"69"),
   372 => (x"0e",x"00",x"0a",x"64"),
   373 => (x"5d",x"5c",x"5b",x"5e"),
   374 => (x"ff",x"c3",x"1e",x"0e"),
   375 => (x"4b",x"d4",x"ff",x"4c"),
   376 => (x"d0",x"ff",x"7b",x"74"),
   377 => (x"c0",x"c8",x"48",x"bf"),
   378 => (x"a6",x"c4",x"98",x"c0"),
   379 => (x"c0",x"02",x"6e",x"58"),
   380 => (x"d0",x"ff",x"87",x"d0"),
   381 => (x"c0",x"c8",x"48",x"bf"),
   382 => (x"a6",x"c4",x"98",x"c0"),
   383 => (x"ff",x"05",x"6e",x"58"),
   384 => (x"d0",x"ff",x"87",x"f0"),
   385 => (x"78",x"c3",x"c4",x"48"),
   386 => (x"66",x"d4",x"7b",x"74"),
   387 => (x"f0",x"ff",x"c0",x"1e"),
   388 => (x"f2",x"1e",x"d8",x"c1"),
   389 => (x"86",x"c8",x"87",x"c5"),
   390 => (x"c0",x"02",x"98",x"70"),
   391 => (x"f3",x"da",x"87",x"cd"),
   392 => (x"87",x"f6",x"e9",x"1e"),
   393 => (x"48",x"c1",x"86",x"c4"),
   394 => (x"74",x"87",x"c4",x"c2"),
   395 => (x"7b",x"fe",x"c3",x"7b"),
   396 => (x"66",x"d8",x"4d",x"c0"),
   397 => (x"4a",x"71",x"49",x"bf"),
   398 => (x"72",x"2a",x"b7",x"d8"),
   399 => (x"70",x"98",x"74",x"48"),
   400 => (x"d0",x"4a",x"71",x"7b"),
   401 => (x"48",x"72",x"2a",x"b7"),
   402 => (x"7b",x"70",x"98",x"74"),
   403 => (x"b7",x"c8",x"4a",x"71"),
   404 => (x"74",x"48",x"72",x"2a"),
   405 => (x"71",x"7b",x"70",x"98"),
   406 => (x"70",x"98",x"74",x"48"),
   407 => (x"48",x"66",x"d8",x"7b"),
   408 => (x"a6",x"dc",x"80",x"c4"),
   409 => (x"c2",x"85",x"c1",x"58"),
   410 => (x"04",x"ad",x"b7",x"c0"),
   411 => (x"74",x"87",x"c3",x"ff"),
   412 => (x"74",x"7b",x"74",x"7b"),
   413 => (x"e0",x"da",x"d8",x"7b"),
   414 => (x"6b",x"7b",x"74",x"49"),
   415 => (x"87",x"c6",x"c0",x"05"),
   416 => (x"ff",x"05",x"89",x"c1"),
   417 => (x"7b",x"74",x"87",x"f3"),
   418 => (x"48",x"bf",x"d0",x"ff"),
   419 => (x"98",x"c0",x"c0",x"c8"),
   420 => (x"6e",x"58",x"a6",x"c4"),
   421 => (x"87",x"d0",x"c0",x"02"),
   422 => (x"48",x"bf",x"d0",x"ff"),
   423 => (x"98",x"c0",x"c0",x"c8"),
   424 => (x"6e",x"58",x"a6",x"c4"),
   425 => (x"87",x"f0",x"ff",x"05"),
   426 => (x"c2",x"48",x"d0",x"ff"),
   427 => (x"26",x"48",x"c0",x"78"),
   428 => (x"57",x"87",x"e0",x"ee"),
   429 => (x"65",x"74",x"69",x"72"),
   430 => (x"69",x"61",x"66",x"20"),
   431 => (x"0a",x"64",x"65",x"6c"),
   432 => (x"5b",x"5e",x"0e",x"00"),
   433 => (x"66",x"d0",x"0e",x"5c"),
   434 => (x"4b",x"66",x"cc",x"4c"),
   435 => (x"ee",x"c5",x"4a",x"c0"),
   436 => (x"ff",x"49",x"df",x"cd"),
   437 => (x"ff",x"c3",x"48",x"d4"),
   438 => (x"48",x"bf",x"70",x"78"),
   439 => (x"05",x"a8",x"fe",x"c3"),
   440 => (x"c1",x"87",x"d8",x"c1"),
   441 => (x"c0",x"48",x"e0",x"e4"),
   442 => (x"ac",x"b7",x"c4",x"78"),
   443 => (x"87",x"dc",x"c0",x"04"),
   444 => (x"70",x"87",x"de",x"ec"),
   445 => (x"c4",x"7b",x"71",x"49"),
   446 => (x"e0",x"e4",x"c1",x"83"),
   447 => (x"80",x"71",x"48",x"bf"),
   448 => (x"58",x"e4",x"e4",x"c1"),
   449 => (x"ac",x"b7",x"8c",x"c4"),
   450 => (x"87",x"e4",x"ff",x"03"),
   451 => (x"06",x"ac",x"b7",x"c0"),
   452 => (x"ff",x"87",x"e5",x"c0"),
   453 => (x"ff",x"c3",x"48",x"d4"),
   454 => (x"49",x"bf",x"70",x"78"),
   455 => (x"c3",x"7b",x"97",x"71"),
   456 => (x"83",x"c1",x"98",x"ff"),
   457 => (x"bf",x"e0",x"e4",x"c1"),
   458 => (x"c1",x"80",x"71",x"48"),
   459 => (x"c1",x"58",x"e4",x"e4"),
   460 => (x"ac",x"b7",x"c0",x"8c"),
   461 => (x"87",x"db",x"ff",x"01"),
   462 => (x"c1",x"4a",x"49",x"c1"),
   463 => (x"d2",x"fe",x"05",x"89"),
   464 => (x"48",x"d4",x"ff",x"87"),
   465 => (x"72",x"78",x"ff",x"c3"),
   466 => (x"87",x"c9",x"ec",x"48"),
   467 => (x"5c",x"5b",x"5e",x"0e"),
   468 => (x"c0",x"c8",x"1e",x"0e"),
   469 => (x"4c",x"c0",x"4b",x"c0"),
   470 => (x"c3",x"48",x"d4",x"ff"),
   471 => (x"d0",x"ff",x"78",x"ff"),
   472 => (x"98",x"73",x"48",x"bf"),
   473 => (x"6e",x"58",x"a6",x"c4"),
   474 => (x"87",x"ce",x"c0",x"02"),
   475 => (x"48",x"bf",x"d0",x"ff"),
   476 => (x"a6",x"c4",x"98",x"73"),
   477 => (x"ff",x"05",x"6e",x"58"),
   478 => (x"d0",x"ff",x"87",x"f2"),
   479 => (x"78",x"c3",x"c4",x"48"),
   480 => (x"c3",x"48",x"d4",x"ff"),
   481 => (x"66",x"d0",x"78",x"ff"),
   482 => (x"f0",x"ff",x"c0",x"1e"),
   483 => (x"ec",x"1e",x"d1",x"c1"),
   484 => (x"86",x"c8",x"87",x"c9"),
   485 => (x"99",x"71",x"49",x"70"),
   486 => (x"87",x"d0",x"c0",x"02"),
   487 => (x"66",x"d4",x"1e",x"71"),
   488 => (x"1e",x"e0",x"df",x"1e"),
   489 => (x"cc",x"87",x"e1",x"e4"),
   490 => (x"87",x"ee",x"c0",x"86"),
   491 => (x"d8",x"1e",x"c0",x"c8"),
   492 => (x"cc",x"fc",x"1e",x"66"),
   493 => (x"70",x"86",x"c8",x"87"),
   494 => (x"bf",x"d0",x"ff",x"4c"),
   495 => (x"c4",x"98",x"73",x"48"),
   496 => (x"02",x"6e",x"58",x"a6"),
   497 => (x"ff",x"87",x"ce",x"c0"),
   498 => (x"73",x"48",x"bf",x"d0"),
   499 => (x"58",x"a6",x"c4",x"98"),
   500 => (x"f2",x"ff",x"05",x"6e"),
   501 => (x"48",x"d0",x"ff",x"87"),
   502 => (x"48",x"74",x"78",x"c2"),
   503 => (x"87",x"f5",x"e9",x"26"),
   504 => (x"64",x"61",x"65",x"52"),
   505 => (x"6d",x"6f",x"63",x"20"),
   506 => (x"64",x"6e",x"61",x"6d"),
   507 => (x"69",x"61",x"66",x"20"),
   508 => (x"20",x"64",x"65",x"6c"),
   509 => (x"25",x"20",x"74",x"61"),
   510 => (x"25",x"28",x"20",x"64"),
   511 => (x"00",x"0a",x"29",x"64"),
   512 => (x"5c",x"5b",x"5e",x"0e"),
   513 => (x"c0",x"1e",x"0e",x"5d"),
   514 => (x"f0",x"ff",x"c0",x"1e"),
   515 => (x"ea",x"1e",x"c9",x"c1"),
   516 => (x"86",x"c8",x"87",x"c9"),
   517 => (x"e4",x"c1",x"1e",x"d2"),
   518 => (x"e4",x"fa",x"1e",x"f2"),
   519 => (x"c0",x"86",x"c8",x"87"),
   520 => (x"d2",x"85",x"c1",x"4d"),
   521 => (x"ff",x"04",x"ad",x"b7"),
   522 => (x"e4",x"c1",x"87",x"f7"),
   523 => (x"49",x"bf",x"97",x"f2"),
   524 => (x"c1",x"99",x"c0",x"c3"),
   525 => (x"c0",x"05",x"a9",x"c0"),
   526 => (x"e4",x"c1",x"87",x"e8"),
   527 => (x"49",x"bf",x"97",x"f9"),
   528 => (x"e4",x"c1",x"31",x"d0"),
   529 => (x"4a",x"bf",x"97",x"fa"),
   530 => (x"b1",x"72",x"32",x"c8"),
   531 => (x"97",x"fb",x"e4",x"c1"),
   532 => (x"b1",x"72",x"4a",x"bf"),
   533 => (x"ff",x"ff",x"ff",x"cf"),
   534 => (x"c1",x"4d",x"71",x"99"),
   535 => (x"c2",x"35",x"ca",x"85"),
   536 => (x"e4",x"c1",x"87",x"ef"),
   537 => (x"4b",x"bf",x"97",x"fb"),
   538 => (x"9b",x"c6",x"33",x"c1"),
   539 => (x"97",x"fc",x"e4",x"c1"),
   540 => (x"b7",x"c7",x"49",x"bf"),
   541 => (x"c1",x"b3",x"71",x"29"),
   542 => (x"bf",x"97",x"f7",x"e4"),
   543 => (x"cf",x"48",x"71",x"49"),
   544 => (x"58",x"a6",x"c4",x"98"),
   545 => (x"97",x"f8",x"e4",x"c1"),
   546 => (x"9c",x"c3",x"4c",x"bf"),
   547 => (x"e4",x"c1",x"34",x"ca"),
   548 => (x"49",x"bf",x"97",x"f9"),
   549 => (x"b4",x"71",x"31",x"c2"),
   550 => (x"97",x"fa",x"e4",x"c1"),
   551 => (x"c0",x"c3",x"49",x"bf"),
   552 => (x"29",x"b7",x"c6",x"99"),
   553 => (x"1e",x"74",x"b4",x"71"),
   554 => (x"73",x"1e",x"66",x"c4"),
   555 => (x"d7",x"e4",x"c0",x"1e"),
   556 => (x"87",x"d4",x"e0",x"1e"),
   557 => (x"83",x"c2",x"86",x"d0"),
   558 => (x"30",x"73",x"48",x"c1"),
   559 => (x"1e",x"73",x"4b",x"70"),
   560 => (x"1e",x"c4",x"e5",x"c0"),
   561 => (x"c8",x"87",x"c1",x"e0"),
   562 => (x"6e",x"48",x"c1",x"86"),
   563 => (x"58",x"a6",x"c4",x"30"),
   564 => (x"81",x"c1",x"49",x"74"),
   565 => (x"b7",x"73",x"4d",x"71"),
   566 => (x"75",x"1e",x"6e",x"95"),
   567 => (x"cd",x"e5",x"c0",x"1e"),
   568 => (x"e3",x"df",x"ff",x"1e"),
   569 => (x"6e",x"86",x"cc",x"87"),
   570 => (x"b7",x"c0",x"c8",x"48"),
   571 => (x"d4",x"c0",x"06",x"a8"),
   572 => (x"6e",x"35",x"c1",x"87"),
   573 => (x"28",x"b7",x"c1",x"48"),
   574 => (x"6e",x"58",x"a6",x"c4"),
   575 => (x"b7",x"c0",x"c8",x"48"),
   576 => (x"ec",x"ff",x"01",x"a8"),
   577 => (x"c0",x"1e",x"75",x"87"),
   578 => (x"ff",x"1e",x"e3",x"e5"),
   579 => (x"c8",x"87",x"f9",x"de"),
   580 => (x"26",x"48",x"75",x"86"),
   581 => (x"63",x"87",x"fc",x"e4"),
   582 => (x"7a",x"69",x"73",x"5f"),
   583 => (x"75",x"6d",x"5f",x"65"),
   584 => (x"20",x"3a",x"74",x"6c"),
   585 => (x"20",x"2c",x"64",x"25"),
   586 => (x"64",x"61",x"65",x"72"),
   587 => (x"5f",x"6c",x"62",x"5f"),
   588 => (x"3a",x"6e",x"65",x"6c"),
   589 => (x"2c",x"64",x"25",x"20"),
   590 => (x"69",x"73",x"63",x"20"),
   591 => (x"20",x"3a",x"65",x"7a"),
   592 => (x"00",x"0a",x"64",x"25"),
   593 => (x"74",x"6c",x"75",x"4d"),
   594 => (x"0a",x"64",x"25",x"20"),
   595 => (x"20",x"64",x"25",x"00"),
   596 => (x"63",x"6f",x"6c",x"62"),
   597 => (x"6f",x"20",x"73",x"6b"),
   598 => (x"69",x"73",x"20",x"66"),
   599 => (x"25",x"20",x"65",x"7a"),
   600 => (x"25",x"00",x"0a",x"64"),
   601 => (x"6c",x"62",x"20",x"64"),
   602 => (x"73",x"6b",x"63",x"6f"),
   603 => (x"20",x"66",x"6f",x"20"),
   604 => (x"20",x"32",x"31",x"35"),
   605 => (x"65",x"74",x"79",x"62"),
   606 => (x"43",x"00",x"0a",x"73"),
   607 => (x"0e",x"00",x"44",x"4d"),
   608 => (x"c0",x"0e",x"5b",x"5e"),
   609 => (x"48",x"66",x"d0",x"4b"),
   610 => (x"06",x"a8",x"b7",x"c0"),
   611 => (x"c8",x"87",x"f6",x"c0"),
   612 => (x"4a",x"bf",x"97",x"66"),
   613 => (x"ba",x"82",x"c0",x"fe"),
   614 => (x"c1",x"48",x"66",x"c8"),
   615 => (x"58",x"a6",x"cc",x"80"),
   616 => (x"bf",x"97",x"66",x"cc"),
   617 => (x"81",x"c0",x"fe",x"49"),
   618 => (x"48",x"66",x"cc",x"b9"),
   619 => (x"a6",x"d0",x"80",x"c1"),
   620 => (x"aa",x"b7",x"71",x"58"),
   621 => (x"c1",x"87",x"c4",x"02"),
   622 => (x"c1",x"87",x"cc",x"48"),
   623 => (x"b7",x"66",x"d0",x"83"),
   624 => (x"ca",x"ff",x"04",x"ab"),
   625 => (x"c4",x"48",x"c0",x"87"),
   626 => (x"26",x"4d",x"26",x"87"),
   627 => (x"26",x"4b",x"26",x"4c"),
   628 => (x"5b",x"5e",x"0e",x"4f"),
   629 => (x"c1",x"0e",x"5d",x"5c"),
   630 => (x"c0",x"48",x"cc",x"ed"),
   631 => (x"e5",x"c1",x"c1",x"78"),
   632 => (x"f5",x"da",x"ff",x"1e"),
   633 => (x"c1",x"86",x"c4",x"87"),
   634 => (x"c0",x"1e",x"c4",x"e5"),
   635 => (x"87",x"dc",x"f5",x"1e"),
   636 => (x"98",x"70",x"86",x"c8"),
   637 => (x"c0",x"87",x"cf",x"05"),
   638 => (x"ff",x"1e",x"d1",x"fe"),
   639 => (x"c4",x"87",x"db",x"da"),
   640 => (x"cb",x"48",x"c0",x"86"),
   641 => (x"c1",x"c1",x"87",x"d6"),
   642 => (x"da",x"ff",x"1e",x"f2"),
   643 => (x"86",x"c4",x"87",x"cc"),
   644 => (x"ed",x"c1",x"4b",x"c0"),
   645 => (x"78",x"c1",x"48",x"f8"),
   646 => (x"c2",x"c1",x"1e",x"c8"),
   647 => (x"e5",x"c1",x"1e",x"c9"),
   648 => (x"da",x"fd",x"1e",x"fa"),
   649 => (x"70",x"86",x"cc",x"87"),
   650 => (x"87",x"c6",x"05",x"98"),
   651 => (x"48",x"f8",x"ed",x"c1"),
   652 => (x"1e",x"c8",x"78",x"c0"),
   653 => (x"1e",x"d2",x"c2",x"c1"),
   654 => (x"1e",x"d6",x"e6",x"c1"),
   655 => (x"cc",x"87",x"c0",x"fd"),
   656 => (x"05",x"98",x"70",x"86"),
   657 => (x"ed",x"c1",x"87",x"c6"),
   658 => (x"78",x"c0",x"48",x"f8"),
   659 => (x"bf",x"f8",x"ed",x"c1"),
   660 => (x"db",x"c2",x"c1",x"1e"),
   661 => (x"ef",x"d9",x"ff",x"1e"),
   662 => (x"c1",x"86",x"c8",x"87"),
   663 => (x"02",x"bf",x"f8",x"ed"),
   664 => (x"c1",x"87",x"d8",x"c2"),
   665 => (x"c1",x"4d",x"c4",x"e5"),
   666 => (x"c1",x"4c",x"c2",x"ec"),
   667 => (x"bf",x"9f",x"c2",x"ed"),
   668 => (x"c1",x"1e",x"71",x"49"),
   669 => (x"c1",x"49",x"c2",x"ed"),
   670 => (x"71",x"89",x"c4",x"e5"),
   671 => (x"c8",x"1e",x"d0",x"1e"),
   672 => (x"ff",x"c0",x"1e",x"c0"),
   673 => (x"d8",x"ff",x"1e",x"c3"),
   674 => (x"86",x"d4",x"87",x"fe"),
   675 => (x"81",x"c8",x"49",x"74"),
   676 => (x"ed",x"c1",x"4b",x"69"),
   677 => (x"49",x"bf",x"9f",x"c2"),
   678 => (x"a9",x"ea",x"d6",x"c5"),
   679 => (x"87",x"d0",x"c0",x"05"),
   680 => (x"81",x"c8",x"49",x"74"),
   681 => (x"d3",x"d9",x"1e",x"69"),
   682 => (x"70",x"86",x"c4",x"87"),
   683 => (x"87",x"df",x"c0",x"4b"),
   684 => (x"fe",x"c7",x"49",x"75"),
   685 => (x"49",x"69",x"9f",x"81"),
   686 => (x"a9",x"d5",x"e9",x"ca"),
   687 => (x"87",x"cf",x"c0",x"02"),
   688 => (x"1e",x"e5",x"fe",x"c0"),
   689 => (x"87",x"d2",x"d7",x"ff"),
   690 => (x"48",x"c0",x"86",x"c4"),
   691 => (x"73",x"87",x"cd",x"c8"),
   692 => (x"c0",x"c0",x"c1",x"1e"),
   693 => (x"ef",x"d7",x"ff",x"1e"),
   694 => (x"c1",x"86",x"c8",x"87"),
   695 => (x"73",x"1e",x"c4",x"e5"),
   696 => (x"87",x"e8",x"f1",x"1e"),
   697 => (x"98",x"70",x"86",x"c8"),
   698 => (x"87",x"c5",x"c0",x"05"),
   699 => (x"eb",x"c7",x"48",x"c0"),
   700 => (x"d8",x"c0",x"c1",x"87"),
   701 => (x"e1",x"d6",x"ff",x"1e"),
   702 => (x"c1",x"86",x"c4",x"87"),
   703 => (x"ff",x"1e",x"ee",x"c2"),
   704 => (x"c4",x"87",x"c5",x"d7"),
   705 => (x"c1",x"1e",x"c8",x"86"),
   706 => (x"c1",x"1e",x"c6",x"c3"),
   707 => (x"f9",x"1e",x"d6",x"e6"),
   708 => (x"86",x"cc",x"87",x"ed"),
   709 => (x"c0",x"05",x"98",x"70"),
   710 => (x"ed",x"c1",x"87",x"c9"),
   711 => (x"78",x"c1",x"48",x"cc"),
   712 => (x"c8",x"87",x"e4",x"c0"),
   713 => (x"cf",x"c3",x"c1",x"1e"),
   714 => (x"fa",x"e5",x"c1",x"1e"),
   715 => (x"87",x"cf",x"f9",x"1e"),
   716 => (x"98",x"70",x"86",x"cc"),
   717 => (x"87",x"cf",x"c0",x"02"),
   718 => (x"1e",x"ff",x"c0",x"c1"),
   719 => (x"87",x"c8",x"d6",x"ff"),
   720 => (x"48",x"c0",x"86",x"c4"),
   721 => (x"c1",x"87",x"d5",x"c6"),
   722 => (x"bf",x"97",x"c2",x"ed"),
   723 => (x"a9",x"d5",x"c1",x"49"),
   724 => (x"87",x"cd",x"c0",x"05"),
   725 => (x"97",x"c3",x"ed",x"c1"),
   726 => (x"ea",x"c2",x"49",x"bf"),
   727 => (x"c5",x"c0",x"02",x"a9"),
   728 => (x"c5",x"48",x"c0",x"87"),
   729 => (x"e5",x"c1",x"87",x"f6"),
   730 => (x"49",x"bf",x"97",x"c4"),
   731 => (x"02",x"a9",x"e9",x"c3"),
   732 => (x"c1",x"87",x"d2",x"c0"),
   733 => (x"bf",x"97",x"c4",x"e5"),
   734 => (x"a9",x"eb",x"c3",x"49"),
   735 => (x"87",x"c5",x"c0",x"02"),
   736 => (x"d7",x"c5",x"48",x"c0"),
   737 => (x"cf",x"e5",x"c1",x"87"),
   738 => (x"71",x"49",x"bf",x"97"),
   739 => (x"cc",x"c0",x"05",x"99"),
   740 => (x"d0",x"e5",x"c1",x"87"),
   741 => (x"c2",x"49",x"bf",x"97"),
   742 => (x"c5",x"c0",x"02",x"a9"),
   743 => (x"c4",x"48",x"c0",x"87"),
   744 => (x"e5",x"c1",x"87",x"fa"),
   745 => (x"48",x"bf",x"97",x"d1"),
   746 => (x"58",x"c8",x"ed",x"c1"),
   747 => (x"bf",x"c4",x"ed",x"c1"),
   748 => (x"c1",x"4a",x"71",x"49"),
   749 => (x"cc",x"ed",x"c1",x"8a"),
   750 => (x"71",x"1e",x"72",x"5a"),
   751 => (x"d8",x"c3",x"c1",x"1e"),
   752 => (x"c3",x"d4",x"ff",x"1e"),
   753 => (x"c1",x"86",x"cc",x"87"),
   754 => (x"bf",x"97",x"d2",x"e5"),
   755 => (x"c1",x"81",x"73",x"49"),
   756 => (x"bf",x"97",x"d3",x"e5"),
   757 => (x"72",x"32",x"c8",x"4a"),
   758 => (x"c1",x"80",x"71",x"48"),
   759 => (x"c1",x"58",x"dc",x"ed"),
   760 => (x"bf",x"97",x"d4",x"e5"),
   761 => (x"f0",x"ed",x"c1",x"48"),
   762 => (x"cc",x"ed",x"c1",x"58"),
   763 => (x"da",x"c2",x"02",x"bf"),
   764 => (x"c1",x"1e",x"c8",x"87"),
   765 => (x"c1",x"1e",x"dc",x"c1"),
   766 => (x"f6",x"1e",x"d6",x"e6"),
   767 => (x"86",x"cc",x"87",x"c1"),
   768 => (x"c0",x"02",x"98",x"70"),
   769 => (x"48",x"c0",x"87",x"c5"),
   770 => (x"c1",x"87",x"d1",x"c3"),
   771 => (x"4a",x"bf",x"c4",x"ed"),
   772 => (x"30",x"c4",x"48",x"72"),
   773 => (x"58",x"f4",x"ed",x"c1"),
   774 => (x"5a",x"ec",x"ed",x"c1"),
   775 => (x"97",x"e9",x"e5",x"c1"),
   776 => (x"31",x"c8",x"49",x"bf"),
   777 => (x"97",x"e8",x"e5",x"c1"),
   778 => (x"81",x"73",x"4b",x"bf"),
   779 => (x"97",x"ea",x"e5",x"c1"),
   780 => (x"33",x"d0",x"4b",x"bf"),
   781 => (x"e5",x"c1",x"81",x"73"),
   782 => (x"4b",x"bf",x"97",x"eb"),
   783 => (x"81",x"73",x"33",x"d8"),
   784 => (x"59",x"f8",x"ed",x"c1"),
   785 => (x"bf",x"ec",x"ed",x"c1"),
   786 => (x"d8",x"ed",x"c1",x"91"),
   787 => (x"ed",x"c1",x"81",x"bf"),
   788 => (x"e5",x"c1",x"59",x"e0"),
   789 => (x"4b",x"bf",x"97",x"f1"),
   790 => (x"e5",x"c1",x"33",x"c8"),
   791 => (x"4c",x"bf",x"97",x"f0"),
   792 => (x"e5",x"c1",x"83",x"74"),
   793 => (x"4c",x"bf",x"97",x"f2"),
   794 => (x"83",x"74",x"34",x"d0"),
   795 => (x"97",x"f3",x"e5",x"c1"),
   796 => (x"9c",x"cf",x"4c",x"bf"),
   797 => (x"83",x"74",x"34",x"d8"),
   798 => (x"5b",x"e4",x"ed",x"c1"),
   799 => (x"92",x"73",x"8b",x"c2"),
   800 => (x"80",x"71",x"48",x"72"),
   801 => (x"58",x"e8",x"ed",x"c1"),
   802 => (x"c1",x"87",x"cf",x"c1"),
   803 => (x"bf",x"97",x"d6",x"e5"),
   804 => (x"c1",x"31",x"c8",x"49"),
   805 => (x"bf",x"97",x"d5",x"e5"),
   806 => (x"c1",x"81",x"72",x"4a"),
   807 => (x"c5",x"59",x"f4",x"ed"),
   808 => (x"81",x"ff",x"c7",x"31"),
   809 => (x"ed",x"c1",x"29",x"c9"),
   810 => (x"e5",x"c1",x"59",x"ec"),
   811 => (x"4a",x"bf",x"97",x"db"),
   812 => (x"e5",x"c1",x"32",x"c8"),
   813 => (x"4b",x"bf",x"97",x"da"),
   814 => (x"ed",x"c1",x"82",x"73"),
   815 => (x"ed",x"c1",x"5a",x"f8"),
   816 => (x"c1",x"92",x"bf",x"ec"),
   817 => (x"82",x"bf",x"d8",x"ed"),
   818 => (x"5a",x"e8",x"ed",x"c1"),
   819 => (x"48",x"e0",x"ed",x"c1"),
   820 => (x"48",x"72",x"78",x"c0"),
   821 => (x"ed",x"c1",x"80",x"71"),
   822 => (x"48",x"c1",x"58",x"e0"),
   823 => (x"0e",x"87",x"ea",x"f3"),
   824 => (x"0e",x"5c",x"5b",x"5e"),
   825 => (x"bf",x"cc",x"ed",x"c1"),
   826 => (x"87",x"cf",x"c0",x"02"),
   827 => (x"c7",x"4a",x"66",x"cc"),
   828 => (x"66",x"cc",x"2a",x"b7"),
   829 => (x"9b",x"ff",x"c1",x"4b"),
   830 => (x"cc",x"87",x"cc",x"c0"),
   831 => (x"b7",x"c8",x"4a",x"66"),
   832 => (x"4b",x"66",x"cc",x"2a"),
   833 => (x"c1",x"9b",x"ff",x"c3"),
   834 => (x"c1",x"1e",x"c4",x"e5"),
   835 => (x"49",x"bf",x"d8",x"ed"),
   836 => (x"1e",x"71",x"81",x"72"),
   837 => (x"c8",x"87",x"f5",x"e8"),
   838 => (x"05",x"98",x"70",x"86"),
   839 => (x"c0",x"87",x"c5",x"c0"),
   840 => (x"87",x"ea",x"c0",x"48"),
   841 => (x"bf",x"cc",x"ed",x"c1"),
   842 => (x"87",x"d4",x"c0",x"02"),
   843 => (x"b7",x"c4",x"49",x"73"),
   844 => (x"c4",x"e5",x"c1",x"91"),
   845 => (x"cf",x"4c",x"69",x"81"),
   846 => (x"ff",x"ff",x"ff",x"ff"),
   847 => (x"87",x"cc",x"c0",x"9c"),
   848 => (x"b7",x"c2",x"49",x"73"),
   849 => (x"c4",x"e5",x"c1",x"91"),
   850 => (x"4c",x"69",x"9f",x"81"),
   851 => (x"fa",x"f1",x"48",x"74"),
   852 => (x"5b",x"5e",x"0e",x"87"),
   853 => (x"f4",x"0e",x"5d",x"5c"),
   854 => (x"76",x"4b",x"c0",x"86"),
   855 => (x"e0",x"ed",x"c1",x"48"),
   856 => (x"80",x"c4",x"78",x"bf"),
   857 => (x"bf",x"e4",x"ed",x"c1"),
   858 => (x"cc",x"ed",x"c1",x"78"),
   859 => (x"ca",x"c0",x"02",x"bf"),
   860 => (x"c4",x"ed",x"c1",x"87"),
   861 => (x"31",x"c4",x"49",x"bf"),
   862 => (x"c1",x"87",x"c7",x"c0"),
   863 => (x"49",x"bf",x"e8",x"ed"),
   864 => (x"a6",x"cc",x"31",x"c4"),
   865 => (x"c8",x"4d",x"c0",x"59"),
   866 => (x"a8",x"c0",x"48",x"66"),
   867 => (x"87",x"f1",x"c2",x"06"),
   868 => (x"99",x"cf",x"49",x"75"),
   869 => (x"87",x"db",x"c0",x"05"),
   870 => (x"1e",x"c4",x"e5",x"c1"),
   871 => (x"48",x"49",x"66",x"c8"),
   872 => (x"a6",x"cc",x"80",x"c1"),
   873 => (x"e6",x"1e",x"71",x"58"),
   874 => (x"86",x"c8",x"87",x"e2"),
   875 => (x"4b",x"c4",x"e5",x"c1"),
   876 => (x"c0",x"87",x"c3",x"c0"),
   877 => (x"6b",x"97",x"83",x"e0"),
   878 => (x"02",x"99",x"71",x"49"),
   879 => (x"97",x"87",x"f9",x"c1"),
   880 => (x"e5",x"c3",x"49",x"6b"),
   881 => (x"ef",x"c1",x"02",x"a9"),
   882 => (x"cb",x"49",x"73",x"87"),
   883 => (x"49",x"69",x"97",x"81"),
   884 => (x"c1",x"05",x"99",x"d8"),
   885 => (x"1e",x"73",x"87",x"e2"),
   886 => (x"87",x"fe",x"ca",x"ff"),
   887 => (x"1e",x"cb",x"86",x"c4"),
   888 => (x"1e",x"66",x"e4",x"c0"),
   889 => (x"d6",x"ee",x"1e",x"73"),
   890 => (x"70",x"86",x"cc",x"87"),
   891 => (x"c7",x"c1",x"05",x"98"),
   892 => (x"dc",x"4a",x"73",x"87"),
   893 => (x"49",x"66",x"dc",x"82"),
   894 => (x"79",x"6a",x"81",x"c4"),
   895 => (x"82",x"da",x"4a",x"73"),
   896 => (x"c8",x"49",x"66",x"dc"),
   897 => (x"48",x"6a",x"9f",x"81"),
   898 => (x"4c",x"71",x"79",x"70"),
   899 => (x"bf",x"cc",x"ed",x"c1"),
   900 => (x"87",x"d2",x"c0",x"02"),
   901 => (x"81",x"d4",x"49",x"73"),
   902 => (x"c0",x"49",x"69",x"9f"),
   903 => (x"71",x"99",x"ff",x"ff"),
   904 => (x"c0",x"32",x"d0",x"4a"),
   905 => (x"4a",x"c0",x"87",x"c2"),
   906 => (x"80",x"6c",x"48",x"72"),
   907 => (x"66",x"dc",x"7c",x"70"),
   908 => (x"c1",x"78",x"c0",x"48"),
   909 => (x"87",x"c0",x"c1",x"48"),
   910 => (x"66",x"c8",x"85",x"c1"),
   911 => (x"cf",x"fd",x"04",x"ad"),
   912 => (x"cc",x"ed",x"c1",x"87"),
   913 => (x"ed",x"c0",x"02",x"bf"),
   914 => (x"fa",x"1e",x"6e",x"87"),
   915 => (x"86",x"c4",x"87",x"d1"),
   916 => (x"6e",x"58",x"a6",x"c4"),
   917 => (x"ff",x"ff",x"cf",x"49"),
   918 => (x"a9",x"99",x"f8",x"ff"),
   919 => (x"87",x"d6",x"c0",x"02"),
   920 => (x"89",x"c2",x"49",x"6e"),
   921 => (x"bf",x"c4",x"ed",x"c1"),
   922 => (x"dc",x"ed",x"c1",x"91"),
   923 => (x"80",x"71",x"48",x"bf"),
   924 => (x"fc",x"58",x"a6",x"c8"),
   925 => (x"48",x"c0",x"87",x"cf"),
   926 => (x"cc",x"ed",x"8e",x"f4"),
   927 => (x"5b",x"5e",x"0e",x"87"),
   928 => (x"bf",x"66",x"c8",x"0e"),
   929 => (x"c8",x"81",x"c1",x"49"),
   930 => (x"09",x"79",x"09",x"66"),
   931 => (x"bf",x"c8",x"ed",x"c1"),
   932 => (x"d0",x"c0",x"05",x"99"),
   933 => (x"4b",x"66",x"c8",x"87"),
   934 => (x"1e",x"6b",x"83",x"c8"),
   935 => (x"c4",x"87",x"c0",x"f9"),
   936 => (x"71",x"49",x"70",x"86"),
   937 => (x"ec",x"48",x"c1",x"7b"),
   938 => (x"5e",x"0e",x"87",x"e3"),
   939 => (x"dc",x"ed",x"c1",x"0e"),
   940 => (x"66",x"c4",x"49",x"bf"),
   941 => (x"6a",x"82",x"c8",x"4a"),
   942 => (x"c1",x"8a",x"c2",x"4a"),
   943 => (x"92",x"bf",x"c4",x"ed"),
   944 => (x"ed",x"c1",x"81",x"72"),
   945 => (x"c4",x"4a",x"bf",x"c8"),
   946 => (x"72",x"9a",x"bf",x"66"),
   947 => (x"1e",x"66",x"c8",x"81"),
   948 => (x"f7",x"e1",x"1e",x"71"),
   949 => (x"70",x"86",x"c8",x"87"),
   950 => (x"c5",x"c0",x"05",x"98"),
   951 => (x"c0",x"48",x"c0",x"87"),
   952 => (x"48",x"c1",x"87",x"c2"),
   953 => (x"0e",x"87",x"e8",x"eb"),
   954 => (x"0e",x"5c",x"5b",x"5e"),
   955 => (x"c1",x"1e",x"66",x"cc"),
   956 => (x"f9",x"1e",x"fc",x"ed"),
   957 => (x"86",x"c8",x"87",x"db"),
   958 => (x"c1",x"02",x"98",x"70"),
   959 => (x"ee",x"c1",x"87",x"d4"),
   960 => (x"c7",x"49",x"bf",x"c0"),
   961 => (x"29",x"c9",x"81",x"ff"),
   962 => (x"4b",x"c0",x"4c",x"71"),
   963 => (x"1e",x"e9",x"fd",x"c0"),
   964 => (x"87",x"c6",x"c6",x"ff"),
   965 => (x"b7",x"c0",x"86",x"c4"),
   966 => (x"c7",x"c1",x"06",x"ac"),
   967 => (x"1e",x"66",x"d0",x"87"),
   968 => (x"1e",x"fc",x"ed",x"c1"),
   969 => (x"c8",x"87",x"c3",x"fe"),
   970 => (x"05",x"98",x"70",x"86"),
   971 => (x"c0",x"87",x"c5",x"c0"),
   972 => (x"87",x"f2",x"c0",x"48"),
   973 => (x"1e",x"fc",x"ed",x"c1"),
   974 => (x"c4",x"87",x"c2",x"fd"),
   975 => (x"48",x"66",x"d0",x"86"),
   976 => (x"d4",x"80",x"c0",x"c8"),
   977 => (x"83",x"c1",x"58",x"a6"),
   978 => (x"04",x"ab",x"b7",x"74"),
   979 => (x"c0",x"87",x"ce",x"ff"),
   980 => (x"66",x"cc",x"87",x"d2"),
   981 => (x"c2",x"fe",x"c0",x"1e"),
   982 => (x"eb",x"c5",x"ff",x"1e"),
   983 => (x"c0",x"86",x"c8",x"87"),
   984 => (x"87",x"c2",x"c0",x"48"),
   985 => (x"e2",x"e9",x"48",x"c1"),
   986 => (x"65",x"70",x"4f",x"87"),
   987 => (x"20",x"64",x"65",x"6e"),
   988 => (x"65",x"6c",x"69",x"66"),
   989 => (x"6f",x"6c",x"20",x"2c"),
   990 => (x"6e",x"69",x"64",x"61"),
   991 => (x"2e",x"2e",x"2e",x"67"),
   992 => (x"61",x"43",x"00",x"0a"),
   993 => (x"20",x"74",x"27",x"6e"),
   994 => (x"6e",x"65",x"70",x"6f"),
   995 => (x"0a",x"73",x"25",x"20"),
   996 => (x"61",x"65",x"52",x"00"),
   997 => (x"66",x"6f",x"20",x"64"),
   998 => (x"52",x"42",x"4d",x"20"),
   999 => (x"69",x"61",x"66",x"20"),
  1000 => (x"0a",x"64",x"65",x"6c"),
  1001 => (x"20",x"6f",x"4e",x"00"),
  1002 => (x"74",x"72",x"61",x"70"),
  1003 => (x"6f",x"69",x"74",x"69"),
  1004 => (x"69",x"73",x"20",x"6e"),
  1005 => (x"74",x"61",x"6e",x"67"),
  1006 => (x"20",x"65",x"72",x"75"),
  1007 => (x"6e",x"75",x"6f",x"66"),
  1008 => (x"4d",x"00",x"0a",x"64"),
  1009 => (x"69",x"73",x"52",x"42"),
  1010 => (x"20",x"3a",x"65",x"7a"),
  1011 => (x"20",x"2c",x"64",x"25"),
  1012 => (x"74",x"72",x"61",x"70"),
  1013 => (x"6f",x"69",x"74",x"69"),
  1014 => (x"7a",x"69",x"73",x"6e"),
  1015 => (x"25",x"20",x"3a",x"65"),
  1016 => (x"6f",x"20",x"2c",x"64"),
  1017 => (x"65",x"73",x"66",x"66"),
  1018 => (x"66",x"6f",x"20",x"74"),
  1019 => (x"67",x"69",x"73",x"20"),
  1020 => (x"64",x"25",x"20",x"3a"),
  1021 => (x"69",x"73",x"20",x"2c"),
  1022 => (x"78",x"30",x"20",x"67"),
  1023 => (x"00",x"0a",x"78",x"25"),
  1024 => (x"64",x"61",x"65",x"52"),
  1025 => (x"20",x"67",x"6e",x"69"),
  1026 => (x"74",x"6f",x"6f",x"62"),
  1027 => (x"63",x"65",x"73",x"20"),
  1028 => (x"20",x"72",x"6f",x"74"),
  1029 => (x"00",x"0a",x"64",x"25"),
  1030 => (x"64",x"61",x"65",x"52"),
  1031 => (x"6f",x"6f",x"62",x"20"),
  1032 => (x"65",x"73",x"20",x"74"),
  1033 => (x"72",x"6f",x"74",x"63"),
  1034 => (x"6f",x"72",x"66",x"20"),
  1035 => (x"69",x"66",x"20",x"6d"),
  1036 => (x"20",x"74",x"73",x"72"),
  1037 => (x"74",x"72",x"61",x"70"),
  1038 => (x"6f",x"69",x"74",x"69"),
  1039 => (x"55",x"00",x"0a",x"6e"),
  1040 => (x"70",x"75",x"73",x"6e"),
  1041 => (x"74",x"72",x"6f",x"70"),
  1042 => (x"70",x"20",x"64",x"65"),
  1043 => (x"69",x"74",x"72",x"61"),
  1044 => (x"6e",x"6f",x"69",x"74"),
  1045 => (x"70",x"79",x"74",x"20"),
  1046 => (x"00",x"0d",x"21",x"65"),
  1047 => (x"33",x"54",x"41",x"46"),
  1048 => (x"20",x"20",x"20",x"32"),
  1049 => (x"61",x"65",x"52",x"00"),
  1050 => (x"67",x"6e",x"69",x"64"),
  1051 => (x"52",x"42",x"4d",x"20"),
  1052 => (x"42",x"4d",x"00",x"0a"),
  1053 => (x"75",x"73",x"20",x"52"),
  1054 => (x"73",x"65",x"63",x"63"),
  1055 => (x"6c",x"75",x"66",x"73"),
  1056 => (x"72",x"20",x"79",x"6c"),
  1057 => (x"0a",x"64",x"61",x"65"),
  1058 => (x"54",x"41",x"46",x"00"),
  1059 => (x"20",x"20",x"36",x"31"),
  1060 => (x"41",x"46",x"00",x"20"),
  1061 => (x"20",x"32",x"33",x"54"),
  1062 => (x"50",x"00",x"20",x"20"),
  1063 => (x"69",x"74",x"72",x"61"),
  1064 => (x"6e",x"6f",x"69",x"74"),
  1065 => (x"6e",x"75",x"6f",x"63"),
  1066 => (x"64",x"25",x"20",x"74"),
  1067 => (x"75",x"48",x"00",x"0a"),
  1068 => (x"6e",x"69",x"74",x"6e"),
  1069 => (x"6f",x"66",x"20",x"67"),
  1070 => (x"69",x"66",x"20",x"72"),
  1071 => (x"79",x"73",x"65",x"6c"),
  1072 => (x"6d",x"65",x"74",x"73"),
  1073 => (x"41",x"46",x"00",x"0a"),
  1074 => (x"20",x"32",x"33",x"54"),
  1075 => (x"46",x"00",x"20",x"20"),
  1076 => (x"36",x"31",x"54",x"41"),
  1077 => (x"00",x"20",x"20",x"20"),
  1078 => (x"73",x"75",x"6c",x"43"),
  1079 => (x"20",x"72",x"65",x"74"),
  1080 => (x"65",x"7a",x"69",x"73"),
  1081 => (x"64",x"25",x"20",x"3a"),
  1082 => (x"6c",x"43",x"20",x"2c"),
  1083 => (x"65",x"74",x"73",x"75"),
  1084 => (x"61",x"6d",x"20",x"72"),
  1085 => (x"20",x"2c",x"6b",x"73"),
  1086 => (x"00",x"0a",x"64",x"25"),
  1087 => (x"c4",x"0e",x"5e",x"0e"),
  1088 => (x"29",x"d8",x"49",x"66"),
  1089 => (x"c4",x"99",x"ff",x"c3"),
  1090 => (x"2a",x"c8",x"4a",x"66"),
  1091 => (x"9a",x"c0",x"fc",x"cf"),
  1092 => (x"66",x"c4",x"b1",x"72"),
  1093 => (x"c0",x"32",x"c8",x"4a"),
  1094 => (x"c0",x"c0",x"f0",x"ff"),
  1095 => (x"c4",x"b1",x"72",x"9a"),
  1096 => (x"32",x"d8",x"4a",x"66"),
  1097 => (x"c0",x"c0",x"c0",x"ff"),
  1098 => (x"b1",x"72",x"9a",x"c0"),
  1099 => (x"87",x"c6",x"48",x"71"),
  1100 => (x"4c",x"26",x"4d",x"26"),
  1101 => (x"4f",x"26",x"4b",x"26"),
  1102 => (x"c4",x"0e",x"5e",x"0e"),
  1103 => (x"2a",x"c8",x"4a",x"66"),
  1104 => (x"cf",x"9a",x"ff",x"c3"),
  1105 => (x"c4",x"9a",x"ff",x"ff"),
  1106 => (x"31",x"c8",x"49",x"66"),
  1107 => (x"99",x"c0",x"fc",x"cf"),
  1108 => (x"ff",x"cf",x"b1",x"72"),
  1109 => (x"48",x"71",x"99",x"ff"),
  1110 => (x"0e",x"87",x"db",x"ff"),
  1111 => (x"66",x"c4",x"0e",x"5e"),
  1112 => (x"cf",x"29",x"d0",x"49"),
  1113 => (x"c4",x"99",x"ff",x"ff"),
  1114 => (x"32",x"d0",x"4a",x"66"),
  1115 => (x"9a",x"c0",x"c0",x"f0"),
  1116 => (x"48",x"71",x"b1",x"72"),
  1117 => (x"00",x"87",x"ff",x"fe"),
  1118 => (x"5e",x"0e",x"4f",x"4f"),
  1119 => (x"e0",x"1e",x"0e",x"5b"),
  1120 => (x"49",x"72",x"4a",x"bf"),
  1121 => (x"99",x"c0",x"e0",x"c0"),
  1122 => (x"87",x"db",x"c2",x"02"),
  1123 => (x"c3",x"9a",x"ff",x"c3"),
  1124 => (x"c9",x"05",x"aa",x"f0"),
  1125 => (x"d6",x"cc",x"c1",x"87"),
  1126 => (x"c1",x"78",x"c1",x"48"),
  1127 => (x"e0",x"c3",x"87",x"fc"),
  1128 => (x"87",x"c9",x"05",x"aa"),
  1129 => (x"48",x"da",x"cc",x"c1"),
  1130 => (x"ed",x"c1",x"78",x"c1"),
  1131 => (x"aa",x"fa",x"c3",x"87"),
  1132 => (x"87",x"e6",x"c1",x"02"),
  1133 => (x"bf",x"da",x"cc",x"c1"),
  1134 => (x"72",x"87",x"c7",x"02"),
  1135 => (x"81",x"c0",x"c2",x"49"),
  1136 => (x"49",x"72",x"87",x"c2"),
  1137 => (x"cc",x"c1",x"4b",x"71"),
  1138 => (x"c0",x"02",x"bf",x"d6"),
  1139 => (x"49",x"73",x"87",x"e2"),
  1140 => (x"b7",x"29",x"b7",x"c4"),
  1141 => (x"de",x"cc",x"c1",x"91"),
  1142 => (x"cf",x"4a",x"73",x"81"),
  1143 => (x"92",x"b7",x"c2",x"9a"),
  1144 => (x"30",x"72",x"48",x"c1"),
  1145 => (x"ba",x"ff",x"4a",x"70"),
  1146 => (x"98",x"69",x"48",x"72"),
  1147 => (x"87",x"de",x"79",x"70"),
  1148 => (x"b7",x"c4",x"49",x"73"),
  1149 => (x"c1",x"91",x"b7",x"29"),
  1150 => (x"73",x"81",x"de",x"cc"),
  1151 => (x"c2",x"9a",x"cf",x"4a"),
  1152 => (x"48",x"c3",x"92",x"b7"),
  1153 => (x"4a",x"70",x"30",x"72"),
  1154 => (x"b0",x"69",x"48",x"72"),
  1155 => (x"cc",x"c1",x"79",x"70"),
  1156 => (x"78",x"c0",x"48",x"da"),
  1157 => (x"48",x"d6",x"cc",x"c1"),
  1158 => (x"bf",x"e0",x"78",x"c0"),
  1159 => (x"c0",x"49",x"72",x"4a"),
  1160 => (x"05",x"99",x"c0",x"e0"),
  1161 => (x"c5",x"87",x"e5",x"fd"),
  1162 => (x"a6",x"c4",x"87",x"cc"),
  1163 => (x"87",x"c4",x"26",x"58"),
  1164 => (x"4c",x"26",x"4d",x"26"),
  1165 => (x"4f",x"26",x"4b",x"26"),
  1166 => (x"c1",x"0e",x"5e",x"0e"),
  1167 => (x"fe",x"1e",x"de",x"cd"),
  1168 => (x"c4",x"87",x"d7",x"f9"),
  1169 => (x"72",x"4a",x"c0",x"86"),
  1170 => (x"91",x"b7",x"c4",x"49"),
  1171 => (x"81",x"de",x"cc",x"c1"),
  1172 => (x"82",x"c1",x"79",x"c0"),
  1173 => (x"04",x"aa",x"b7",x"d0"),
  1174 => (x"c4",x"87",x"ec",x"ff"),
  1175 => (x"d5",x"ff",x"87",x"e7"),
  1176 => (x"0e",x"5e",x"0e",x"87"),
  1177 => (x"c4",x"49",x"66",x"c4"),
  1178 => (x"91",x"b7",x"29",x"b7"),
  1179 => (x"81",x"de",x"cc",x"c1"),
  1180 => (x"cf",x"4a",x"66",x"c4"),
  1181 => (x"92",x"b7",x"c2",x"9a"),
  1182 => (x"30",x"72",x"48",x"c2"),
  1183 => (x"ba",x"ff",x"4a",x"70"),
  1184 => (x"98",x"69",x"48",x"72"),
  1185 => (x"ed",x"fe",x"79",x"70"),
  1186 => (x"5b",x"5e",x"0e",x"87"),
  1187 => (x"4a",x"66",x"c8",x"0e"),
  1188 => (x"b7",x"2a",x"b7",x"c4"),
  1189 => (x"de",x"cc",x"c1",x"92"),
  1190 => (x"4b",x"66",x"c8",x"82"),
  1191 => (x"b7",x"c2",x"9b",x"cf"),
  1192 => (x"73",x"49",x"6a",x"93"),
  1193 => (x"c2",x"99",x"c3",x"29"),
  1194 => (x"70",x"30",x"73",x"48"),
  1195 => (x"73",x"bb",x"ff",x"4b"),
  1196 => (x"70",x"98",x"6a",x"48"),
  1197 => (x"fd",x"48",x"71",x"7a"),
  1198 => (x"5e",x"0e",x"87",x"fa"),
  1199 => (x"66",x"c8",x"0e",x"5b"),
  1200 => (x"2a",x"b7",x"c4",x"4a"),
  1201 => (x"cc",x"c1",x"92",x"b7"),
  1202 => (x"66",x"c8",x"82",x"de"),
  1203 => (x"c2",x"99",x"cf",x"49"),
  1204 => (x"48",x"6a",x"91",x"b7"),
  1205 => (x"49",x"70",x"28",x"71"),
  1206 => (x"9b",x"c3",x"4b",x"71"),
  1207 => (x"c0",x"05",x"ab",x"c2"),
  1208 => (x"66",x"c8",x"87",x"e2"),
  1209 => (x"29",x"b7",x"c4",x"49"),
  1210 => (x"cc",x"c1",x"91",x"b7"),
  1211 => (x"66",x"c8",x"81",x"de"),
  1212 => (x"c2",x"9a",x"cf",x"4a"),
  1213 => (x"48",x"c2",x"92",x"b7"),
  1214 => (x"4a",x"70",x"30",x"72"),
  1215 => (x"48",x"72",x"ba",x"ff"),
  1216 => (x"79",x"70",x"98",x"69"),
  1217 => (x"c0",x"02",x"ab",x"c2"),
  1218 => (x"49",x"c0",x"87",x"c5"),
  1219 => (x"c1",x"87",x"c2",x"c0"),
  1220 => (x"fc",x"48",x"71",x"49"),
  1221 => (x"00",x"00",x"87",x"de"),
  1222 => (x"00",x"00",x"00",x"00"),
  1223 => (x"00",x"00",x"00",x"00"),
  1224 => (x"06",x"06",x"00",x"00"),
  1225 => (x"06",x"06",x"06",x"06"),
  1226 => (x"06",x"06",x"06",x"06"),
  1227 => (x"06",x"06",x"06",x"06"),
  1228 => (x"06",x"06",x"06",x"06"),
  1229 => (x"06",x"06",x"06",x"06"),
  1230 => (x"06",x"06",x"06",x"06"),
  1231 => (x"06",x"06",x"06",x"06"),
  1232 => (x"06",x"06",x"06",x"06"),
  1233 => (x"06",x"06",x"06",x"06"),
  1234 => (x"06",x"06",x"06",x"06"),
  1235 => (x"06",x"06",x"06",x"06"),
  1236 => (x"06",x"06",x"06",x"06"),
  1237 => (x"06",x"06",x"06",x"06"),
  1238 => (x"06",x"06",x"06",x"06"),
  1239 => (x"65",x"4b",x"06",x"06"),
  1240 => (x"61",x"6f",x"62",x"79"),
  1241 => (x"69",x"20",x"64",x"72"),
  1242 => (x"20",x"74",x"69",x"6e"),
  1243 => (x"63",x"6e",x"75",x"66"),
  1244 => (x"6e",x"6f",x"69",x"74"),
  1245 => (x"fe",x"1e",x"00",x"0a"),
  1246 => (x"c6",x"48",x"bf",x"f0"),
  1247 => (x"26",x"4d",x"26",x"87"),
  1248 => (x"26",x"4b",x"26",x"4c"),
  1249 => (x"f0",x"fe",x"1e",x"4f"),
  1250 => (x"f6",x"78",x"c1",x"48"),
  1251 => (x"f0",x"fe",x"1e",x"87"),
  1252 => (x"ee",x"78",x"c0",x"48"),
  1253 => (x"0e",x"5e",x"0e",x"87"),
  1254 => (x"bf",x"e0",x"d3",x"c1"),
  1255 => (x"c1",x"31",x"cb",x"49"),
  1256 => (x"4a",x"bf",x"dc",x"d3"),
  1257 => (x"b1",x"72",x"32",x"c8"),
  1258 => (x"87",x"c6",x"48",x"71"),
  1259 => (x"4c",x"26",x"4d",x"26"),
  1260 => (x"4f",x"26",x"4b",x"26"),
  1261 => (x"48",x"c0",x"f8",x"1e"),
  1262 => (x"c1",x"78",x"66",x"c4"),
  1263 => (x"c0",x"48",x"d4",x"d3"),
  1264 => (x"1e",x"87",x"ef",x"78"),
  1265 => (x"48",x"d8",x"d3",x"c1"),
  1266 => (x"d3",x"c1",x"78",x"c0"),
  1267 => (x"66",x"c4",x"48",x"d4"),
  1268 => (x"c5",x"1e",x"c0",x"78"),
  1269 => (x"ff",x"86",x"c4",x"87"),
  1270 => (x"5e",x"0e",x"87",x"d8"),
  1271 => (x"0e",x"5d",x"5c",x"5b"),
  1272 => (x"ff",x"c0",x"4a",x"c0"),
  1273 => (x"48",x"66",x"d0",x"4d"),
  1274 => (x"bf",x"d8",x"d3",x"c1"),
  1275 => (x"d9",x"c1",x"02",x"a8"),
  1276 => (x"49",x"66",x"d0",x"87"),
  1277 => (x"cb",x"02",x"99",x"c1"),
  1278 => (x"d4",x"d3",x"c1",x"87"),
  1279 => (x"88",x"c1",x"48",x"bf"),
  1280 => (x"58",x"d8",x"d3",x"c1"),
  1281 => (x"c2",x"49",x"66",x"d0"),
  1282 => (x"87",x"cb",x"02",x"99"),
  1283 => (x"bf",x"d4",x"d3",x"c1"),
  1284 => (x"c1",x"80",x"c1",x"48"),
  1285 => (x"c1",x"58",x"d8",x"d3"),
  1286 => (x"48",x"bf",x"d4",x"d3"),
  1287 => (x"03",x"a8",x"b7",x"c0"),
  1288 => (x"d3",x"c1",x"87",x"c6"),
  1289 => (x"78",x"c1",x"48",x"d4"),
  1290 => (x"bf",x"d4",x"d3",x"c1"),
  1291 => (x"a8",x"b7",x"c1",x"48"),
  1292 => (x"c1",x"87",x"c6",x"06"),
  1293 => (x"c0",x"48",x"d4",x"d3"),
  1294 => (x"49",x"66",x"d0",x"78"),
  1295 => (x"c2",x"02",x"99",x"d0"),
  1296 => (x"c1",x"4a",x"c1",x"87"),
  1297 => (x"d0",x"48",x"d8",x"d3"),
  1298 => (x"d3",x"c1",x"78",x"66"),
  1299 => (x"c0",x"49",x"bf",x"d4"),
  1300 => (x"87",x"c8",x"02",x"a9"),
  1301 => (x"d7",x"02",x"a9",x"c1"),
  1302 => (x"87",x"eb",x"c0",x"87"),
  1303 => (x"bf",x"dc",x"d3",x"c1"),
  1304 => (x"c3",x"81",x"72",x"49"),
  1305 => (x"e0",x"d3",x"c1",x"99"),
  1306 => (x"c5",x"4b",x"71",x"59"),
  1307 => (x"87",x"df",x"93",x"b7"),
  1308 => (x"d3",x"c1",x"4b",x"d4"),
  1309 => (x"72",x"49",x"bf",x"e0"),
  1310 => (x"e4",x"d3",x"c1",x"b9"),
  1311 => (x"05",x"99",x"71",x"59"),
  1312 => (x"4d",x"d7",x"87",x"cd"),
  1313 => (x"c1",x"87",x"c8",x"c0"),
  1314 => (x"4b",x"bf",x"d4",x"d3"),
  1315 => (x"f8",x"93",x"b7",x"c5"),
  1316 => (x"0d",x"7d",x"0d",x"c4"),
  1317 => (x"c0",x"93",x"b7",x"c3"),
  1318 => (x"e6",x"d3",x"c1",x"4c"),
  1319 => (x"97",x"82",x"73",x"4a"),
  1320 => (x"32",x"d0",x"4a",x"6a"),
  1321 => (x"49",x"e5",x"d3",x"c1"),
  1322 => (x"69",x"97",x"81",x"73"),
  1323 => (x"71",x"31",x"c8",x"49"),
  1324 => (x"e4",x"d3",x"c1",x"b2"),
  1325 => (x"97",x"81",x"73",x"49"),
  1326 => (x"b2",x"71",x"49",x"69"),
  1327 => (x"b7",x"c4",x"49",x"74"),
  1328 => (x"81",x"c8",x"f8",x"91"),
  1329 => (x"83",x"c3",x"79",x"72"),
  1330 => (x"b7",x"c5",x"84",x"c1"),
  1331 => (x"c8",x"ff",x"04",x"ac"),
  1332 => (x"87",x"d8",x"fb",x"87"),
  1333 => (x"00",x"00",x"00",x"00"),
  1334 => (x"00",x"00",x"00",x"00"),
  1335 => (x"00",x"00",x"00",x"03"),
  1336 => (x"00",x"00",x"00",x"00"),
  1337 => (x"55",x"00",x"3b",x"db"),
  1338 => (x"49",x"d5",x"00",x"48"),
  1339 => (x"00",x"48",x"51",x"00"),
  1340 => (x"cf",x"00",x"3b",x"d1"),
  1341 => (x"05",x"21",x"08",x"b8"),
  1342 => (x"02",x"19",x"27",x"05"),
  1343 => (x"2f",x"02",x"21",x"e1"),
  1344 => (x"9c",x"c9",x"02",x"1d"),
  1345 => (x"04",x"a5",x"29",x"03"),
  1346 => (x"e9",x"04",x"a5",x"2f"),
  1347 => (x"a5",x"29",x"04",x"9d"),
  1348 => (x"07",x"bc",x"ef",x"03"),
  1349 => (x"27",x"00",x"85",x"21"),
  1350 => (x"84",x"e1",x"03",x"9d"),
  1351 => (x"07",x"bd",x"21",x"00"),
  1352 => (x"29",x"fb",x"3d",x"26"),
  1353 => (x"9d",x"e1",x"24",x"85"),
  1354 => (x"27",x"85",x"29",x"24"),
  1355 => (x"61",x"24",x"bd",x"26"),
  1356 => (x"52",x"91",x"01",x"cc"),
  1357 => (x"02",x"52",x"91",x"02"),
  1358 => (x"67",x"02",x"5e",x"91"),
  1359 => (x"1c",x"ef",x"a9",x"d2"),
  1360 => (x"94",x"a5",x"21",x"73"),
  1361 => (x"e1",x"94",x"a5",x"27"),
  1362 => (x"25",x"2f",x"74",x"9c"),
  1363 => (x"5b",x"5e",x"0e",x"93"),
  1364 => (x"f8",x"0e",x"5d",x"5c"),
  1365 => (x"c0",x"48",x"76",x"86"),
  1366 => (x"f7",x"e3",x"c1",x"78"),
  1367 => (x"f9",x"ec",x"fe",x"1e"),
  1368 => (x"fe",x"86",x"c4",x"87"),
  1369 => (x"70",x"87",x"f0",x"fd"),
  1370 => (x"87",x"cd",x"02",x"98"),
  1371 => (x"87",x"e1",x"d1",x"ff"),
  1372 => (x"c4",x"02",x"98",x"70"),
  1373 => (x"c2",x"49",x"c1",x"87"),
  1374 => (x"71",x"49",x"c0",x"87"),
  1375 => (x"f0",x"c2",x"02",x"99"),
  1376 => (x"cd",x"e4",x"c1",x"87"),
  1377 => (x"c8",x"ee",x"c1",x"1e"),
  1378 => (x"c4",x"df",x"ff",x"1e"),
  1379 => (x"70",x"86",x"c8",x"87"),
  1380 => (x"dc",x"c2",x"02",x"98"),
  1381 => (x"48",x"a6",x"c4",x"87"),
  1382 => (x"bf",x"cc",x"ee",x"c1"),
  1383 => (x"f8",x"1e",x"c1",x"78"),
  1384 => (x"86",x"c4",x"87",x"d2"),
  1385 => (x"da",x"f8",x"1e",x"c5"),
  1386 => (x"c1",x"86",x"c4",x"87"),
  1387 => (x"fe",x"1e",x"fa",x"e2"),
  1388 => (x"c4",x"87",x"e7",x"eb"),
  1389 => (x"c1",x"48",x"f8",x"86"),
  1390 => (x"02",x"66",x"c4",x"78"),
  1391 => (x"c4",x"87",x"db",x"c1"),
  1392 => (x"e5",x"c1",x"4c",x"66"),
  1393 => (x"ee",x"c1",x"1e",x"c4"),
  1394 => (x"dd",x"e3",x"1e",x"c8"),
  1395 => (x"70",x"86",x"c8",x"87"),
  1396 => (x"87",x"c5",x"05",x"98"),
  1397 => (x"d7",x"cb",x"48",x"c0"),
  1398 => (x"b7",x"c0",x"c8",x"87"),
  1399 => (x"87",x"c6",x"04",x"ac"),
  1400 => (x"8c",x"4a",x"c0",x"c8"),
  1401 => (x"4a",x"74",x"87",x"c4"),
  1402 => (x"e5",x"c1",x"4c",x"c0"),
  1403 => (x"49",x"72",x"4b",x"c4"),
  1404 => (x"99",x"71",x"8a",x"c1"),
  1405 => (x"13",x"87",x"d4",x"02"),
  1406 => (x"80",x"c0",x"fe",x"48"),
  1407 => (x"78",x"08",x"fc",x"b8"),
  1408 => (x"c1",x"49",x"72",x"08"),
  1409 => (x"05",x"99",x"71",x"8a"),
  1410 => (x"c1",x"87",x"ec",x"ff"),
  1411 => (x"e1",x"1e",x"c8",x"ee"),
  1412 => (x"86",x"c4",x"87",x"eb"),
  1413 => (x"fe",x"05",x"9c",x"74"),
  1414 => (x"48",x"f8",x"87",x"e8"),
  1415 => (x"e3",x"c1",x"78",x"c0"),
  1416 => (x"e9",x"fe",x"1e",x"d3"),
  1417 => (x"86",x"c4",x"87",x"f4"),
  1418 => (x"c7",x"f6",x"1e",x"c0"),
  1419 => (x"de",x"86",x"c4",x"87"),
  1420 => (x"f5",x"1e",x"c1",x"87"),
  1421 => (x"86",x"c4",x"87",x"fe"),
  1422 => (x"c6",x"f6",x"1e",x"c6"),
  1423 => (x"c1",x"86",x"c4",x"87"),
  1424 => (x"fe",x"1e",x"d9",x"e3"),
  1425 => (x"c4",x"87",x"d3",x"e9"),
  1426 => (x"87",x"eb",x"ec",x"86"),
  1427 => (x"c0",x"87",x"fa",x"ff"),
  1428 => (x"48",x"a6",x"c4",x"4b"),
  1429 => (x"4d",x"4c",x"78",x"c0"),
  1430 => (x"f0",x"1e",x"d8",x"c1"),
  1431 => (x"86",x"c4",x"87",x"eb"),
  1432 => (x"c0",x"02",x"98",x"70"),
  1433 => (x"e0",x"c0",x"87",x"c3"),
  1434 => (x"f0",x"1e",x"d2",x"b4"),
  1435 => (x"86",x"c4",x"87",x"db"),
  1436 => (x"c0",x"02",x"98",x"70"),
  1437 => (x"b4",x"d0",x"87",x"c2"),
  1438 => (x"cc",x"f0",x"1e",x"d4"),
  1439 => (x"70",x"86",x"c4",x"87"),
  1440 => (x"c3",x"c0",x"02",x"98"),
  1441 => (x"b4",x"e0",x"c0",x"87"),
  1442 => (x"fc",x"ef",x"1e",x"d1"),
  1443 => (x"70",x"86",x"c4",x"87"),
  1444 => (x"c2",x"c0",x"02",x"98"),
  1445 => (x"dd",x"b4",x"d0",x"87"),
  1446 => (x"87",x"ed",x"ef",x"1e"),
  1447 => (x"98",x"70",x"86",x"c4"),
  1448 => (x"87",x"c2",x"c0",x"02"),
  1449 => (x"1e",x"db",x"b4",x"c1"),
  1450 => (x"c4",x"87",x"de",x"ef"),
  1451 => (x"02",x"98",x"70",x"86"),
  1452 => (x"c2",x"87",x"c2",x"c0"),
  1453 => (x"ef",x"1e",x"dc",x"b4"),
  1454 => (x"86",x"c4",x"87",x"cf"),
  1455 => (x"c0",x"02",x"98",x"70"),
  1456 => (x"b4",x"c4",x"87",x"c2"),
  1457 => (x"ee",x"1e",x"e3",x"c0"),
  1458 => (x"86",x"c4",x"87",x"ff"),
  1459 => (x"c0",x"02",x"98",x"70"),
  1460 => (x"b4",x"c8",x"87",x"c2"),
  1461 => (x"ee",x"1e",x"da",x"c1"),
  1462 => (x"86",x"c4",x"87",x"ef"),
  1463 => (x"c0",x"02",x"98",x"70"),
  1464 => (x"b3",x"d0",x"87",x"c2"),
  1465 => (x"ee",x"1e",x"d9",x"c1"),
  1466 => (x"86",x"c4",x"87",x"df"),
  1467 => (x"c0",x"02",x"98",x"70"),
  1468 => (x"e0",x"c0",x"87",x"c3"),
  1469 => (x"1e",x"d4",x"c2",x"b3"),
  1470 => (x"c4",x"87",x"ce",x"ee"),
  1471 => (x"02",x"98",x"70",x"86"),
  1472 => (x"d0",x"87",x"c2",x"c0"),
  1473 => (x"1e",x"d1",x"c2",x"b3"),
  1474 => (x"c4",x"87",x"fe",x"ed"),
  1475 => (x"02",x"98",x"70",x"86"),
  1476 => (x"c0",x"87",x"c3",x"c0"),
  1477 => (x"f5",x"c3",x"b3",x"e0"),
  1478 => (x"87",x"ed",x"ed",x"1e"),
  1479 => (x"98",x"70",x"86",x"c4"),
  1480 => (x"87",x"c2",x"c0",x"02"),
  1481 => (x"f2",x"c3",x"b3",x"c1"),
  1482 => (x"87",x"dd",x"ed",x"1e"),
  1483 => (x"98",x"70",x"86",x"c4"),
  1484 => (x"87",x"c2",x"c0",x"02"),
  1485 => (x"eb",x"c3",x"b3",x"c2"),
  1486 => (x"87",x"cd",x"ed",x"1e"),
  1487 => (x"98",x"70",x"86",x"c4"),
  1488 => (x"87",x"c2",x"c0",x"02"),
  1489 => (x"f4",x"c3",x"b3",x"c4"),
  1490 => (x"87",x"fd",x"ec",x"1e"),
  1491 => (x"98",x"70",x"86",x"c4"),
  1492 => (x"87",x"c2",x"c0",x"02"),
  1493 => (x"f1",x"c0",x"b3",x"c8"),
  1494 => (x"87",x"ed",x"ec",x"1e"),
  1495 => (x"98",x"70",x"86",x"c4"),
  1496 => (x"87",x"c8",x"c0",x"02"),
  1497 => (x"d0",x"48",x"66",x"c4"),
  1498 => (x"58",x"a6",x"c8",x"b0"),
  1499 => (x"ec",x"1e",x"f2",x"c0"),
  1500 => (x"86",x"c4",x"87",x"d7"),
  1501 => (x"c0",x"02",x"98",x"70"),
  1502 => (x"66",x"c4",x"87",x"c9"),
  1503 => (x"b0",x"e0",x"c0",x"48"),
  1504 => (x"c1",x"58",x"a6",x"c8"),
  1505 => (x"c0",x"ec",x"1e",x"c3"),
  1506 => (x"70",x"86",x"c4",x"87"),
  1507 => (x"c8",x"c0",x"02",x"98"),
  1508 => (x"48",x"66",x"c4",x"87"),
  1509 => (x"a6",x"c8",x"b0",x"c1"),
  1510 => (x"1e",x"c2",x"c1",x"58"),
  1511 => (x"c4",x"87",x"ea",x"eb"),
  1512 => (x"02",x"98",x"70",x"86"),
  1513 => (x"c4",x"87",x"c8",x"c0"),
  1514 => (x"b0",x"c2",x"48",x"66"),
  1515 => (x"c0",x"58",x"a6",x"c8"),
  1516 => (x"d4",x"eb",x"1e",x"fb"),
  1517 => (x"70",x"86",x"c4",x"87"),
  1518 => (x"c8",x"c0",x"02",x"98"),
  1519 => (x"48",x"66",x"c4",x"87"),
  1520 => (x"a6",x"c8",x"b0",x"c4"),
  1521 => (x"1e",x"cb",x"c1",x"58"),
  1522 => (x"c4",x"87",x"fe",x"ea"),
  1523 => (x"02",x"98",x"70",x"86"),
  1524 => (x"c4",x"87",x"c8",x"c0"),
  1525 => (x"b0",x"c8",x"48",x"66"),
  1526 => (x"c0",x"58",x"a6",x"c8"),
  1527 => (x"e8",x"ea",x"1e",x"ee"),
  1528 => (x"70",x"86",x"c4",x"87"),
  1529 => (x"c2",x"c0",x"02",x"98"),
  1530 => (x"c0",x"b5",x"c1",x"87"),
  1531 => (x"d8",x"ea",x"1e",x"f6"),
  1532 => (x"70",x"86",x"c4",x"87"),
  1533 => (x"c2",x"c0",x"02",x"98"),
  1534 => (x"c0",x"b5",x"c2",x"87"),
  1535 => (x"c8",x"ea",x"1e",x"fd"),
  1536 => (x"70",x"86",x"c4",x"87"),
  1537 => (x"c2",x"c0",x"02",x"98"),
  1538 => (x"d6",x"b5",x"c4",x"87"),
  1539 => (x"87",x"f9",x"e9",x"1e"),
  1540 => (x"98",x"70",x"86",x"c4"),
  1541 => (x"87",x"c2",x"c0",x"02"),
  1542 => (x"1e",x"de",x"b5",x"c8"),
  1543 => (x"c4",x"87",x"ea",x"e9"),
  1544 => (x"02",x"98",x"70",x"86"),
  1545 => (x"d0",x"87",x"c2",x"c0"),
  1546 => (x"1e",x"e6",x"c0",x"b5"),
  1547 => (x"c4",x"87",x"da",x"e9"),
  1548 => (x"02",x"98",x"70",x"86"),
  1549 => (x"c0",x"87",x"c3",x"c0"),
  1550 => (x"1e",x"c7",x"b5",x"e0"),
  1551 => (x"c4",x"87",x"fb",x"e9"),
  1552 => (x"02",x"98",x"70",x"86"),
  1553 => (x"c7",x"87",x"fb",x"c0"),
  1554 => (x"87",x"d5",x"e8",x"1e"),
  1555 => (x"48",x"6e",x"86",x"c4"),
  1556 => (x"a6",x"c4",x"b8",x"c1"),
  1557 => (x"ed",x"1e",x"6e",x"58"),
  1558 => (x"86",x"c4",x"87",x"da"),
  1559 => (x"e3",x"c1",x"1e",x"6e"),
  1560 => (x"e1",x"fe",x"1e",x"e9"),
  1561 => (x"86",x"c8",x"87",x"e2"),
  1562 => (x"d5",x"c0",x"05",x"6e"),
  1563 => (x"87",x"e5",x"ec",x"87"),
  1564 => (x"4a",x"71",x"49",x"70"),
  1565 => (x"0a",x"f4",x"b2",x"c1"),
  1566 => (x"0a",x"f4",x"0a",x"7a"),
  1567 => (x"09",x"f4",x"0a",x"7a"),
  1568 => (x"c4",x"fd",x"09",x"79"),
  1569 => (x"73",x"0d",x"7d",x"0d"),
  1570 => (x"c4",x"31",x"d0",x"49"),
  1571 => (x"32",x"c8",x"4a",x"66"),
  1572 => (x"48",x"71",x"b1",x"72"),
  1573 => (x"c8",x"fd",x"b0",x"74"),
  1574 => (x"6e",x"08",x"78",x"08"),
  1575 => (x"87",x"c7",x"c0",x"02"),
  1576 => (x"f5",x"ec",x"1e",x"73"),
  1577 => (x"e3",x"86",x"c4",x"87"),
  1578 => (x"cd",x"e3",x"87",x"cd"),
  1579 => (x"87",x"df",x"f6",x"87"),
  1580 => (x"4d",x"26",x"8e",x"f8"),
  1581 => (x"4b",x"26",x"4c",x"26"),
  1582 => (x"70",x"4f",x"4f",x"26"),
  1583 => (x"64",x"65",x"6e",x"65"),
  1584 => (x"6c",x"69",x"66",x"20"),
  1585 => (x"6c",x"20",x"2c",x"65"),
  1586 => (x"69",x"64",x"61",x"6f"),
  1587 => (x"2e",x"2e",x"67",x"6e"),
  1588 => (x"44",x"00",x"0a",x"2e"),
  1589 => (x"0a",x"65",x"6e",x"6f"),
  1590 => (x"20",x"44",x"53",x"00"),
  1591 => (x"74",x"6f",x"6f",x"62"),
  1592 => (x"69",x"61",x"66",x"20"),
  1593 => (x"0a",x"64",x"65",x"6c"),
  1594 => (x"6f",x"68",x"53",x"00"),
  1595 => (x"65",x"6d",x"20",x"77"),
  1596 => (x"25",x"20",x"75",x"6e"),
  1597 => (x"49",x"00",x"0a",x"64"),
  1598 => (x"69",x"74",x"69",x"6e"),
  1599 => (x"7a",x"69",x"6c",x"61"),
  1600 => (x"20",x"67",x"6e",x"69"),
  1601 => (x"63",x"20",x"44",x"53"),
  1602 => (x"0a",x"64",x"72",x"61"),
  1603 => (x"4d",x"41",x"52",x"00"),
  1604 => (x"45",x"47",x"41",x"50"),
  1605 => (x"4d",x"4f",x"52",x"20"),
  1606 => (x"00",x"12",x"38",x"00"),
  1607 => (x"00",x"12",x"38",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
